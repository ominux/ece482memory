* # FILE NAME: /HOME/ENGR/TRUTY1/CADENCE/SIMULATION/WHOLE_CKT/HSPICES/          
* SCHEMATIC/NETLIST/WHOLE_CKT.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON NOV 16 12:59:16 2009
   
* GLOBAL NET DEFINITIONS
.lib "/apps/Linux/cadence-Sept2009/ncsu-cdk-1.5.1/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "/apps/Linux/cadence-Sept2009/ncsu-cdk-1.5.1/models/hspice/public/publicModel/tsmc18dN" NMOS 

.GLOBAL VDD! 
* FILE NAME: ECE482MEMORY_WHOLE_CKT_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: WHOLE_CKT.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
XI62 A0 A1 A2 CLK DFF_OUT_6 DFF_OUT_5 DFF_OUT_4 DFF_OUT_3 DFF_OUT_2 DFF_OUT_1 
+DFF_OUT_0 H_3 H_2 H_1 H_0 OUT_3 OUT_2 OUT_1 OUT_0 _DFF_OUT_6 _DFF_OUT_5 
+_DFF_OUT_4 _DFF_OUT_3 _DFF_OUT_2 _DFF_OUT_1 _DFF_OUT_0 0 VDD! PART1_G1 
C0 OUT_3 0  50E-15 M=1.0 
C3 OUT_0 0  50E-15 M=1.0 
C2 OUT_1 0  50E-15 M=1.0 
C1 OUT_2 0  50E-15 M=1.0 
XI52 CLK CLK_D2__ INV_1 
XI59 CLK_D3_ CLK_D3 INV_2 
XI56 CLK_D1__ NET066 INV_3 
XI58 CLK_D2 CLK_D2_ INV_4 
XI49 CLK CLK_D1_ INV_5 
XI54 NET067 CLK_D3_ INV_4 
XI61 NET068 NET067 INV_5 
XI53 CLK NET068 INV_6 
XI39 CLK CLK_D0_ INV_7 
XI50 NET066 CLK_D1 INV_8 
XI51 CLK_D2__ CLK_D2 INV_9 
XI55 CLK_D1_ CLK_D1__ INV_3 
VA2_GEN A2 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 6.4E-9 12.8E-9 
V1 CLK 0  PULSE 0.0 1.8 0.0 80E-12 80E-12 700E-12 1.6E-9 
VA0_GEN A0 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 1.6E-9 3.2E-9 
VA1_GEN A1 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 3.2E-9 6.4E-9 
V0 VDD! 0  1.8 
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_7 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(450E-9) AD=+2.02500000E-13 
+AS=+2.02500000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(900E-9) AD=+4.05000000E-13 
+AS=+4.05000000E-13 PD=+2.70000000E-06 PS=+2.70000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_7 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_6 A Y 
M0 Y A 0 0  TSMC18DN  L=(270E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(270E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_6 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_4 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(810E-9) AD=+3.64500000E-13 
+AS=+3.64500000E-13 PD=+2.52000000E-06 PS=+2.52000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_4 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_3 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_3 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(1.08E-6) AD=+4.86000000E-13 
+AS=+4.86000000E-13 PD=+3.06000000E-06 PS=+3.06000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_8 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_8 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_9 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(720E-9) AD=+3.24000000E-13 
+AS=+3.24000000E-13 PD=+2.34000000E-06 PS=+2.34000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_9 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:43 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_5 A Y 
M0 Y A 0 0  TSMC18DN  L=(270E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(270E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_5 
   
   
   
* FILE NAME: ECE482MEMORY_PART1_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: PART1.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 15:31:42 2009.
   
* TERMINAL MAPPING: A0 = A0
*                   A1 = A1
*                   A2 = A2
*                   CLK = CLK
*                   DFF_OUT<6> = DFF_OUT_6
*                   DFF_OUT<5> = DFF_OUT_5
*                   DFF_OUT<4> = DFF_OUT_4
*                   DFF_OUT<3> = DFF_OUT_3
*                   DFF_OUT<2> = DFF_OUT_2
*                   DFF_OUT<1> = DFF_OUT_1
*                   DFF_OUT<0> = DFF_OUT_0
*                   H<3> = H_3
*                   H<2> = H_2
*                   H<1> = H_1
*                   H<0> = H_0
*                   OUT<3> = OUT_3
*                   OUT<2> = OUT_2
*                   OUT<1> = OUT_1
*                   OUT<0> = OUT_0
*                   _DFF_OUT<6> = _DFF_OUT_6
*                   _DFF_OUT<5> = _DFF_OUT_5
*                   _DFF_OUT<4> = _DFF_OUT_4
*                   _DFF_OUT<3> = _DFF_OUT_3
*                   _DFF_OUT<2> = _DFF_OUT_2
*                   _DFF_OUT<1> = _DFF_OUT_1
*                   _DFF_OUT<0> = _DFF_OUT_0
*                   GND = GND
*                   VDD = VDD
.SUBCKT PART1_G1 A0 A1 A2 CLK DFF_OUT_6 DFF_OUT_5 DFF_OUT_4 DFF_OUT_3 
+DFF_OUT_2 DFF_OUT_1 DFF_OUT_0 H_3 H_2 H_1 H_0 OUT_3 OUT_2 OUT_1 OUT_0 
+_DFF_OUT_6 _DFF_OUT_5 _DFF_OUT_4 _DFF_OUT_3 _DFF_OUT_2 _DFF_OUT_1 _DFF_OUT_0 
+GND VDD 
C190 VDD 143  38.4992999999998E-18 M=1.0 
C191 VDD 139  51.8561999999999E-18 M=1.0 
C192 VDD 128  58.1418E-18 M=1.0 
C193 VDD 102  26.7138000000001E-18 M=1.0 
C194 VDD _DFF_OUT_4  58.1418E-18 M=1.0 
C195 _DFF_OUT_2 VDD  40.0707E-18 M=1.0 
C196 GND 143  58.9275000000002E-18 M=1.0 
C197 GND 119  32.2137E-18 M=1.0 
C198 GND 118  32.2137E-18 M=1.0 
C199 GND 117  32.2137E-18 M=1.0 
C200 GND 116  32.2137E-18 M=1.0 
C201 GND 115  32.2137000000001E-18 M=1.0 
C202 GND 114  32.2137E-18 M=1.0 
C203 GND 113  32.2137000000001E-18 M=1.0 
C204 GND 102  109.998E-18 M=1.0 
C205 GND 95  39.285E-18 M=1.0 
C206 GND 16  230.9958E-18 M=1.0 
C207 GND _DFF_OUT_4  201.9249E-18 M=1.0 
C208 GND _DFF_OUT_3  206.6391E-18 M=1.0 
C209 GND _DFF_OUT_2  149.283E-18 M=1.0 
C210 CLK GND  206.6391E-18 M=1.0 
C211 _DFF_OUT_0 GND  206.6391E-18 M=1.0 
C212 DFF_OUT_4 GND  36.1422000000002E-18 M=1.0 
C213 _DFF_OUT_6 VDD  40.0707E-18 M=1.0 
C214 _DFF_OUT_6 GND  149.283E-18 M=1.0 
C215 112 114  62.3646E-18 M=1.0 
C216 102 111  62.3646E-18 M=1.0 
C217 95 112  62.3646E-18 M=1.0 
C218 95 111  62.3646E-18 M=1.0 
C219 67 84  62.3646E-18 M=1.0 
C220 67 76  62.3646E-18 M=1.0 
C221 67 70  62.3646E-18 M=1.0 
C222 60 70  62.3646E-18 M=1.0 
C223 28 74  62.3646E-18 M=1.0 
C224 26 84  62.3646E-18 M=1.0 
C225 16 74  62.3646E-18 M=1.0 
C226 1 81  62.3646E-18 M=1.0 
C227 1 10  62.3646E-18 M=1.0 
C228 VDD 143  46.3662000000001E-18 M=1.0 
C229 VDD 120  57.3146999999998E-18 M=1.0 
C230 VDD 118  56.6991E-18 M=1.0 
C231 VDD 116  56.6991E-18 M=1.0 
C232 VDD 114  56.6991E-18 M=1.0 
C233 VDD 102  54.2808E-18 M=1.0 
C234 VDD 95  56.6991E-18 M=1.0 
C235 VDD 88  79.0029E-18 M=1.0 
C236 VDD 81  99.0584999999999E-18 M=1.0 
C237 VDD 10  99.0584999999998E-18 M=1.0 
C238 VDD DFF_OUT_1  54.2808E-18 M=1.0 
C239 _DFF_OUT_3 VDD  27.1404E-18 M=1.0 
C240 DFF_OUT_0 VDD  27.1404E-18 M=1.0 
C241 _DFF_OUT_2 DFF_OUT_0  62.3646E-18 M=1.0 
C242 _DFF_OUT_1 VDD  27.1404E-18 M=1.0 
C243 GND 133  448.4826E-18 M=1.0 
C244 GND 124  94.068E-18 M=1.0 
C245 GND 119  209.3463E-18 M=1.0 
C246 GND 116  209.3463E-18 M=1.0 
C247 GND 115  209.3463E-18 M=1.0 
C248 GND 114  209.3463E-18 M=1.0 
C249 GND 111  314.4501E-18 M=1.0 
C250 GND 102  176.4513E-18 M=1.0 
C251 GND 95  195.0066E-18 M=1.0 
C252 GND 88  203.13E-18 M=1.0 
C253 GND 81  163.881E-18 M=1.0 
C254 GND 10  163.881E-18 M=1.0 
C255 GND 3  442.1286E-18 M=1.0 
C256 GND DFF_OUT_1  467.829000000001E-18 M=1.0 
C257 GND DFF_OUT_0  1.0597635E-15 M=1.0 
C258 CLK VDD  187.9047E-18 M=1.0 
C259 CLK GND  204.3828E-18 M=1.0 
C260 _DFF_OUT_0 VDD  27.1404E-18 M=1.0 
C261 _DFF_OUT_0 GND  170.2845E-18 M=1.0 
C262 _DFF_OUT_6 VDD  176.8356E-18 M=1.0 
C263 _DFF_OUT_6 DFF_OUT_4  152.442E-18 M=1.0 
C264 DFF_OUT_2 _DFF_OUT_0  62.3646E-18 M=1.0 
C265 112 114  55.3986E-18 M=1.0 
C266 102 111  104.8338E-18 M=1.0 
C267 95 111  119.3148E-18 M=1.0 
C268 95 102  297.5607E-18 M=1.0 
C269 81 110  55.3986E-18 M=1.0 
C270 67 93  65.0448E-18 M=1.0 
C271 67 84  65.0448E-18 M=1.0 
C272 67 76  65.0448E-18 M=1.0 
C273 67 70  65.0448E-18 M=1.0 
C274 60 76  65.0448E-18 M=1.0 
C275 60 70  65.0448E-18 M=1.0 
C276 28 74  65.0448E-18 M=1.0 
C277 26 93  65.0448E-18 M=1.0 
C278 26 84  65.0448E-18 M=1.0 
C279 23 28  65.0448E-18 M=1.0 
C280 16 74  64.945575E-18 M=1.0 
C281 16 21  65.0448E-18 M=1.0 
C282 10 110  55.3986E-18 M=1.0 
C283 2 74  60.31485E-18 M=1.0 
C284 2 17  60.31485E-18 M=1.0 
C285 1 81  120.3381E-18 M=1.0 
C286 1 10  120.70665E-18 M=1.0 
C287 _DFF_OUT_4 117  299.4885E-18 M=1.0 
C288 VDD 119  34.9776E-18 M=1.0 
C289 VDD 118  34.9776E-18 M=1.0 
C290 VDD 117  34.9776E-18 M=1.0 
C291 VDD 116  34.9776E-18 M=1.0 
C292 VDD 115  34.9776E-18 M=1.0 
C293 VDD 114  34.9776E-18 M=1.0 
C294 VDD 113  34.9776E-18 M=1.0 
C295 VDD 88  55.3986E-18 M=1.0 
C296 VDD 10  65.0448E-18 M=1.0 
C297 _DFF_OUT_3 116  299.4885E-18 M=1.0 
C298 _DFF_OUT_3 VDD  65.5065E-18 M=1.0 
C299 _DFF_OUT_2 115  299.4885E-18 M=1.0 
C300 _DFF_OUT_2 VDD  710.9973E-18 M=1.0 
C301 _DFF_OUT_1 114  299.4885E-18 M=1.0 
C302 _DFF_OUT_1 DFF_OUT_1  111.933E-18 M=1.0 
C303 _DFF_OUT_1 VDD  65.5065E-18 M=1.0 
C304 GND 119  48.9483E-18 M=1.0 
C305 GND 118  48.9483E-18 M=1.0 
C306 GND 117  48.9483E-18 M=1.0 
C307 GND 116  48.9483E-18 M=1.0 
C308 GND 115  48.9483E-18 M=1.0 
C309 GND 114  48.9483E-18 M=1.0 
C310 GND 113  48.9483E-18 M=1.0 
C311 GND 102  157.7223E-18 M=1.0 
C312 GND 95  107.1702E-18 M=1.0 
C313 GND 76  4.232592E-15 M=1.0 
C314 GND 70  3.3164172E-15 M=1.0 
C315 GND 28  2.4578964E-15 M=1.0 
C316 GND 3  23.74515E-18 M=1.0 
C317 GND _DFF_OUT_3  1.3545225E-15 M=1.0 
C318 GND DFF_OUT_0  55.3986E-18 M=1.0 
C319 GND _DFF_OUT_2  4.2521103E-15 M=1.0 
C320 GND _DFF_OUT_1  537.4107E-18 M=1.0 
C321 _DFF_OUT_0 113  299.4885E-18 M=1.0 
C322 _DFF_OUT_0 _DFF_OUT_2  55.3986E-18 M=1.0 
C323 _DFF_OUT_0 GND  2.73641355E-15 M=1.0 
C324 DFF_OUT_6 _DFF_OUT_4  37.944E-18 M=1.0 
C325 DFF_OUT_4 _DFF_OUT_4  55.3986E-18 M=1.0 
C326 DFF_OUT_4 _DFF_OUT_3  55.3986E-18 M=1.0 
C327 DFF_OUT_4 _DFF_OUT_0  69.534E-18 M=1.0 
C328 _DFF_OUT_6 119  299.4885E-18 M=1.0 
C329 _DFF_OUT_6 VDD  327.7071E-18 M=1.0 
C330 _DFF_OUT_6 DFF_OUT_0  55.3986E-18 M=1.0 
C331 _DFF_OUT_6 GND  4.345002E-15 M=1.0 
C332 _DFF_OUT_6 _DFF_OUT_0  55.3986E-18 M=1.0 
C333 DFF_OUT_3 _DFF_OUT_4  110.7972E-18 M=1.0 
C334 _DFF_OUT_5 118  299.4885E-18 M=1.0 
C335 _DFF_OUT_5 DFF_OUT_5  55.3986E-18 M=1.0 
C336 DFF_OUT_2 _DFF_OUT_2  55.3986E-18 M=1.0 
C337 DFF_OUT_2 _DFF_OUT_0  69.3378E-18 M=1.0 
C338 102 112  52.3044E-18 M=1.0 
C339 95 111  37.6677E-18 M=1.0 
C340 3 110  175.510125E-18 M=1.0 
C341 3 93  104.6088E-18 M=1.0 
C342 3 88  37.6677E-18 M=1.0 
C343 3 84  104.6088E-18 M=1.0 
C344 3 81  150.907725E-18 M=1.0 
C345 3 76  104.6088E-18 M=1.0 
C346 3 70  104.6088E-18 M=1.0 
C347 3 28  104.6088E-18 M=1.0 
C348 3 16  104.6088E-18 M=1.0 
C349 3 10  163.433925E-18 M=1.0 
C350 2 3  104.6088E-18 M=1.0 
C351 1 3  104.6088E-18 M=1.0 
C352 VDD 3  388.04715E-18 M=1.0 
C353 _DFF_OUT_2 DFF_OUT_0  173.054925E-18 M=1.0 
C354 _DFF_OUT_1 _DFF_OUT_2  781.97805E-18 M=1.0 
C355 GND 139  200.52585E-18 M=1.0 
C356 GND 3  1.0969011E-15 M=1.0 
C357 GND _DFF_OUT_3  123.4143E-18 M=1.0 
C358 _DFF_OUT_0 _DFF_OUT_1  116.5779E-18 M=1.0 
C359 _DFF_OUT_0 GND  123.4143E-18 M=1.0 
C360 _DFF_OUT_6 _DFF_OUT_2  52.3044E-18 M=1.0 
C361 _DFF_OUT_6 _DFF_OUT_1  52.3044E-18 M=1.0 
C362 DFF_OUT_2 _DFF_OUT_6  52.3044E-18 M=1.0 
C363 DFF_OUT_1 133  495.25155E-18 M=1.0 
C364 _DFF_OUT_2 DFF_OUT_1  49.5477E-18 M=1.0 
C365 _DFF_OUT_6 DFF_OUT_1  49.5477E-18 M=1.0 
C366 VDD 111  362.600549999999E-18 M=1.0 
C367 VDD 110  280.494900000001E-18 M=1.0 
C368 VDD 105  26.7138E-18 M=1.0 
C369 GND 105  109.998E-18 M=1.0 
C370 GND 98  39.285E-18 M=1.0 
C371 GND 84  318.9942E-18 M=1.0 
C372 GND 70  324.4941E-18 M=1.0 
C373 GND 1  230.9958E-18 M=1.0 
C374 GND VDD  958.161150000001E-18 M=1.0 
C375 112 117  62.3646E-18 M=1.0 
C376 105 111  62.3646E-18 M=1.0 
C377 98 112  62.3646E-18 M=1.0 
C378 98 111  62.3646E-18 M=1.0 
C379 73 84  62.3646E-18 M=1.0 
C380 73 76  62.3646E-18 M=1.0 
C381 68 93  62.3646E-18 M=1.0 
C382 68 84  62.3646E-18 M=1.0 
C383 68 76  62.3646E-18 M=1.0 
C384 68 70  62.3646E-18 M=1.0 
C385 1 83  62.3646E-18 M=1.0 
C386 1 82  62.3646E-18 M=1.0 
C387 VDD 117  56.6991E-18 M=1.0 
C388 VDD 110  646.6122E-18 M=1.0 
C389 VDD 105  54.2808E-18 M=1.0 
C390 VDD 98  56.6991E-18 M=1.0 
C391 VDD 89  106.7094E-18 M=1.0 
C392 VDD 83  89.3960999999999E-18 M=1.0 
C393 VDD 82  89.3961000000001E-18 M=1.0 
C394 VDD 5  74.331E-18 M=1.0 
C395 GND 117  209.3463E-18 M=1.0 
C396 GND 105  176.4513E-18 M=1.0 
C397 GND 98  195.0066E-18 M=1.0 
C398 GND 93  478.3374E-18 M=1.0 
C399 GND 90  883.9386E-18 M=1.0 
C400 GND 83  164.9034E-18 M=1.0 
C401 GND 82  164.9034E-18 M=1.0 
C402 GND 1  741.3435E-18 M=1.0 
C403 112 117  55.3986E-18 M=1.0 
C404 105 112  78.3504E-18 M=1.0 
C405 105 111  104.8338E-18 M=1.0 
C406 98 112  50.39325E-18 M=1.0 
C407 98 111  119.3148E-18 M=1.0 
C408 98 105  297.5607E-18 M=1.0 
C409 83 110  55.3986E-18 M=1.0 
C410 82 110  55.3986E-18 M=1.0 
C411 68 93  65.0448E-18 M=1.0 
C412 68 84  65.0448E-18 M=1.0 
C413 68 76  65.0448E-18 M=1.0 
C414 28 68  65.0448E-18 M=1.0 
C415 16 77  60.31485E-18 M=1.0 
C416 2 79  60.31485E-18 M=1.0 
C417 1 110  582.5736E-18 M=1.0 
C418 1 83  55.62945E-18 M=1.0 
C419 1 82  120.3381E-18 M=1.0 
C420 VDD 28  1.6542396E-15 M=1.0 
C421 VDD 16  874.9422E-18 M=1.0 
C422 VDD 5  76.4973E-18 M=1.0 
C423 GND 105  157.7223E-18 M=1.0 
C424 GND 98  107.1702E-18 M=1.0 
C425 GND 83  293.6736E-18 M=1.0 
C426 GND 82  293.6736E-18 M=1.0 
C427 105 112  52.3044E-18 M=1.0 
C428 98 111  37.6677E-18 M=1.0 
C429 5 110  156.9132E-18 M=1.0 
C430 5 90  37.6677E-18 M=1.0 
C431 5 84  104.6088E-18 M=1.0 
C432 5 83  148.216275E-18 M=1.0 
C433 5 28  104.6088E-18 M=1.0 
C434 5 16  104.6088E-18 M=1.0 
C435 4 110  156.9132E-18 M=1.0 
C436 4 93  104.6088E-18 M=1.0 
C437 4 89  37.6677E-18 M=1.0 
C438 4 82  99.2826E-18 M=1.0 
C439 4 28  138.312E-18 M=1.0 
C440 2 5  104.6088E-18 M=1.0 
C441 GND 110  326.0655E-18 M=1.0 
C442 GND 93  230.9958E-18 M=1.0 
C443 GND 76  230.9958E-18 M=1.0 
C444 GND 28  318.9942E-18 M=1.0 
C445 GND 2  307.9944E-18 M=1.0 
C446 58 76  62.3646E-18 M=1.0 
C447 57 76  62.3646E-18 M=1.0 
C448 57 70  62.3646E-18 M=1.0 
C449 25 93  62.3646E-18 M=1.0 
C450 24 93  62.3646E-18 M=1.0 
C451 19 28  62.3646E-18 M=1.0 
C452 16 19  62.3646E-18 M=1.0 
C453 16 18  62.3646E-18 M=1.0 
C454 1 13  62.3646E-18 M=1.0 
C455 1 12  62.3646E-18 M=1.0 
C456 1 11  62.3646E-18 M=1.0 
C457 VDD 13  99.0585E-18 M=1.0 
C458 VDD 12  89.3960999999999E-18 M=1.0 
C459 VDD 11  89.3961000000001E-18 M=1.0 
C460 VDD 4  72.4293E-18 M=1.0 
C461 GND 84  442.683E-18 M=1.0 
C462 GND 70  231.26985E-18 M=1.0 
C463 GND 16  601.947900000001E-18 M=1.0 
C464 GND 13  163.881E-18 M=1.0 
C465 GND 12  164.9034E-18 M=1.0 
C466 GND 11  164.9034E-18 M=1.0 
C467 GND 6  1.5927561E-15 M=1.0 
C468 GND 5  647.3034E-18 M=1.0 
C469 GND 4  254.1132E-18 M=1.0 
C470 68 70  65.0448E-18 M=1.0 
C471 63 70  65.0448E-18 M=1.0 
C472 62 70  65.0448E-18 M=1.0 
C473 61 76  65.0448E-18 M=1.0 
C474 59 84  65.0448E-18 M=1.0 
C475 58 84  65.0448E-18 M=1.0 
C476 58 76  65.0448E-18 M=1.0 
C477 57 84  65.0448E-18 M=1.0 
C478 57 76  65.0448E-18 M=1.0 
C479 57 70  65.0448E-18 M=1.0 
C480 27 93  65.0448E-18 M=1.0 
C481 25 93  65.0448E-18 M=1.0 
C482 25 28  65.0448E-18 M=1.0 
C483 24 93  65.0448E-18 M=1.0 
C484 24 28  65.0448E-18 M=1.0 
C485 19 28  65.0448E-18 M=1.0 
C486 16 22  65.0448E-18 M=1.0 
C487 16 19  65.0448E-18 M=1.0 
C488 16 18  65.0448E-18 M=1.0 
C489 13 110  55.3986E-18 M=1.0 
C490 12 110  55.3986E-18 M=1.0 
C491 11 110  55.3986E-18 M=1.0 
C492 2 20  60.31485E-18 M=1.0 
C493 2 19  60.31485E-18 M=1.0 
C494 2 18  60.31485E-18 M=1.0 
C495 1 13  64.84635E-18 M=1.0 
C496 1 12  120.70665E-18 M=1.0 
C497 1 11  120.70665E-18 M=1.0 
C498 VDD 110  1.3851225E-15 M=1.0 
C499 VDD 84  260.1792E-18 M=1.0 
C500 VDD 76  260.1792E-18 M=1.0 
C501 VDD 70  195.1344E-18 M=1.0 
C502 VDD 13  65.0448E-18 M=1.0 
C503 VDD 12  65.0448E-18 M=1.0 
C504 VDD 11  65.0448E-18 M=1.0 
C505 VDD 2  874.9422E-18 M=1.0 
C506 GND 110  5.6929644E-15 M=1.0 
C507 GND 2  3.4484679E-15 M=1.0 
C508 GND 1  3.1785741E-15 M=1.0 
C509 5 93  104.6088E-18 M=1.0 
C510 5 76  104.6088E-18 M=1.0 
C511 5 70  104.6088E-18 M=1.0 
C512 5 12  161.071875E-18 M=1.0 
C513 4 84  138.312E-18 M=1.0 
C514 4 76  104.6088E-18 M=1.0 
C515 4 70  138.312E-18 M=1.0 
C516 4 16  104.6088E-18 M=1.0 
C517 4 11  113.6682E-18 M=1.0 
C518 2 4  104.6088E-18 M=1.0 
C519 1 5  104.6088E-18 M=1.0 
C520 1 4  104.6088E-18 M=1.0 
C521 VDD 5  185.822325E-18 M=1.0 
C522 VDD 4  134.736975E-18 M=1.0 
C523 GND 5  985.361175E-18 M=1.0 
C524 GND 4  973.752075000001E-18 M=1.0 
C525 VDD 112  252.9954E-18 M=1.0 
C526 VDD 107  26.7138E-18 M=1.0 
C527 VDD 106  26.7138E-18 M=1.0 
C528 GND 111  288.74475E-18 M=1.0 
C529 GND 107  109.998E-18 M=1.0 
C530 GND 106  109.998E-18 M=1.0 
C531 GND 100  39.285E-18 M=1.0 
C532 GND 99  39.285E-18 M=1.0 
C533 112 119  62.3646E-18 M=1.0 
C534 112 118  62.3646E-18 M=1.0 
C535 107 111  62.3646E-18 M=1.0 
C536 106 111  62.3646E-18 M=1.0 
C537 100 112  62.3646E-18 M=1.0 
C538 100 111  62.3646E-18 M=1.0 
C539 99 112  62.3646E-18 M=1.0 
C540 99 111  62.3646E-18 M=1.0 
C541 VDD 119  56.6991E-18 M=1.0 
C542 VDD 111  182.6118E-18 M=1.0 
C543 VDD 107  54.2808E-18 M=1.0 
C544 VDD 106  54.2808E-18 M=1.0 
C545 VDD 100  56.6991E-18 M=1.0 
C546 VDD 99  56.6991E-18 M=1.0 
C547 VDD 90  81.4212E-18 M=1.0 
C548 VDD 6  81.4212E-18 M=1.0 
C549 GND 118  209.3463E-18 M=1.0 
C550 GND 107  176.4513E-18 M=1.0 
C551 GND 106  176.4513E-18 M=1.0 
C552 GND 100  195.0066E-18 M=1.0 
C553 GND 99  195.0066E-18 M=1.0 
C554 112 119  55.3986E-18 M=1.0 
C555 112 118  55.3986E-18 M=1.0 
C556 107 112  78.3504E-18 M=1.0 
C557 107 111  104.8338E-18 M=1.0 
C558 106 112  78.3504E-18 M=1.0 
C559 106 111  104.8338E-18 M=1.0 
C560 100 112  50.39325E-18 M=1.0 
C561 100 111  119.3148E-18 M=1.0 
C562 100 107  297.5607E-18 M=1.0 
C563 99 112  50.39325E-18 M=1.0 
C564 99 111  119.3148E-18 M=1.0 
C565 99 106  297.5607E-18 M=1.0 
C566 VDD 107  65.5065E-18 M=1.0 
C567 VDD 106  65.5065E-18 M=1.0 
C568 VDD 105  65.5065E-18 M=1.0 
C569 VDD 100  34.9776E-18 M=1.0 
C570 VDD 99  34.9776E-18 M=1.0 
C571 VDD 98  34.9776E-18 M=1.0 
C572 VDD 90  55.3986E-18 M=1.0 
C573 VDD 6  55.3986E-18 M=1.0 
C574 GND 112  7.38479385000001E-15 M=1.0 
C575 GND 111  2.95639245E-15 M=1.0 
C576 GND 107  157.7223E-18 M=1.0 
C577 GND 106  157.7223E-18 M=1.0 
C578 GND 100  107.1702E-18 M=1.0 
C579 GND 99  107.1702E-18 M=1.0 
C580 111 112  1.8995076E-15 M=1.0 
C581 106 112  52.3044E-18 M=1.0 
C582 100 111  37.6677E-18 M=1.0 
C583 99 111  37.6677E-18 M=1.0 
C584 VDD 112  1.6100667E-15 M=1.0 
C585 VDD 111  2.24015535E-15 M=1.0 
C586 VDD 104  26.7138E-18 M=1.0 
C587 VDD 103  26.7138E-18 M=1.0 
C588 GND 112  302.4945E-18 M=1.0 
C589 GND 104  109.998E-18 M=1.0 
C590 GND 103  109.998E-18 M=1.0 
C591 GND 97  39.285E-18 M=1.0 
C592 GND 96  39.285E-18 M=1.0 
C593 112 116  62.3646E-18 M=1.0 
C594 112 115  62.3646E-18 M=1.0 
C595 104 111  62.3646E-18 M=1.0 
C596 103 111  62.3646E-18 M=1.0 
C597 97 112  62.3646E-18 M=1.0 
C598 97 111  62.3646E-18 M=1.0 
C599 96 112  62.3646E-18 M=1.0 
C600 96 111  62.3646E-18 M=1.0 
C601 VDD 115  56.6991E-18 M=1.0 
C602 VDD 104  54.2808E-18 M=1.0 
C603 VDD 103  54.2808E-18 M=1.0 
C604 VDD 97  56.6991E-18 M=1.0 
C605 VDD 96  56.6991E-18 M=1.0 
C606 GND 112  377.2269E-18 M=1.0 
C607 GND 104  176.4513E-18 M=1.0 
C608 GND 103  176.4513E-18 M=1.0 
C609 GND 97  195.0066E-18 M=1.0 
C610 GND 96  195.0066E-18 M=1.0 
C611 GND 89  460.3761E-18 M=1.0 
C612 GND VDD  6.01515495E-15 M=1.0 
C613 112 116  55.3986E-18 M=1.0 
C614 112 115  55.3986E-18 M=1.0 
C615 104 112  78.3504E-18 M=1.0 
C616 104 111  104.8338E-18 M=1.0 
C617 103 112  78.3504E-18 M=1.0 
C618 103 111  104.8338E-18 M=1.0 
C619 102 112  78.3504E-18 M=1.0 
C620 97 112  50.39325E-18 M=1.0 
C621 97 111  119.3148E-18 M=1.0 
C622 97 104  297.5607E-18 M=1.0 
C623 96 112  50.39325E-18 M=1.0 
C624 96 111  119.3148E-18 M=1.0 
C625 96 103  297.5607E-18 M=1.0 
C626 95 112  50.39325E-18 M=1.0 
C627 VDD 104  65.5065E-18 M=1.0 
C628 VDD 103  65.5065E-18 M=1.0 
C629 VDD 97  34.9776E-18 M=1.0 
C630 VDD 96  34.9776E-18 M=1.0 
C631 VDD 89  55.3986E-18 M=1.0 
C632 VDD 4  73.85085E-18 M=1.0 
C633 GND 104  157.7223E-18 M=1.0 
C634 GND 103  157.7223E-18 M=1.0 
C635 GND 97  107.1702E-18 M=1.0 
C636 GND 96  107.1702E-18 M=1.0 
C637 104 112  52.3044E-18 M=1.0 
C638 103 112  52.3044E-18 M=1.0 
C639 97 111  37.6677E-18 M=1.0 
C640 96 111  37.6677E-18 M=1.0 
C641 VDD 87  53.4276E-18 M=1.0 
C642 VDD 66  53.4276E-18 M=1.0 
C643 VDD 65  139.0689E-18 M=1.0 
C644 VDD 64  53.4276000000002E-18 M=1.0 
C645 VDD 8  157.925700000001E-18 M=1.0 
C646 GND 108  129.640499999998E-18 M=1.0 
C647 GND 86  369.279000000001E-18 M=1.0 
C648 GND 72  29.8566000000003E-18 M=1.0 
C649 GND 71  29.8566000000001E-18 M=1.0 
C650 GND 64  182.2824E-18 M=1.0 
C651 84 86  62.3646E-18 M=1.0 
C652 76 87  124.7292E-18 M=1.0 
C653 72 108  62.3646E-18 M=1.0 
C654 71 108  62.3646000000001E-18 M=1.0 
C655 70 86  124.7292E-18 M=1.0 
C656 66 84  124.7292E-18 M=1.0 
C657 65 76  62.3646E-18 M=1.0 
C658 65 70  62.3646E-18 M=1.0 
C659 VDD 109  114.8382E-18 M=1.0 
C660 VDD 87  27.1404E-18 M=1.0 
C661 VDD 84  76.0680000000001E-18 M=1.0 
C662 VDD 76  76.0680000000001E-18 M=1.0 
C663 VDD 72  46.674E-18 M=1.0 
C664 VDD 71  46.6740000000001E-18 M=1.0 
C665 VDD 70  76.0680000000001E-18 M=1.0 
C666 VDD 66  61.8380999999999E-18 M=1.0 
C667 VDD 64  54.2808000000002E-18 M=1.0 
C668 VDD 8  59.6339999999999E-18 M=1.0 
C669 VDD A1  27.1404000000001E-18 M=1.0 
C670 GND 110  1.4370291E-15 M=1.0 
C671 GND 109  143.2593E-18 M=1.0 
C672 GND 87  1.2551877E-15 M=1.0 
C673 GND 76  349.0218E-18 M=1.0 
C674 GND 72  205.6968E-18 M=1.0 
C675 GND 71  188.6859E-18 M=1.0 
C676 GND 66  1.4018382E-15 M=1.0 
C677 GND 65  767.791799999999E-18 M=1.0 
C678 GND 64  167.6628E-18 M=1.0 
C679 GND 9  771.4521E-18 M=1.0 
C680 GND A1  65.1743999999999E-18 M=1.0 
C681 CLK 71  62.3646000000001E-18 M=1.0 
C682 CLK 64  62.3646E-18 M=1.0 
C683 86 87  395.226E-18 M=1.0 
C684 84 93  110.7972E-18 M=1.0 
C685 84 86  146.0529E-18 M=1.0 
C686 76 93  110.7972E-18 M=1.0 
C687 76 84  110.7972E-18 M=1.0 
C688 72 108  55.3986E-18 M=1.0 
C689 71 108  75.29535E-18 M=1.0 
C690 70 93  55.3986E-18 M=1.0 
C691 70 84  55.3986E-18 M=1.0 
C692 70 76  55.3986E-18 M=1.0 
C693 66 87  55.3986E-18 M=1.0 
C694 66 86  55.3986E-18 M=1.0 
C695 66 84  55.3986E-18 M=1.0 
C696 66 76  55.3986E-18 M=1.0 
C697 66 70  55.3986E-18 M=1.0 
C698 65 87  221.5944E-18 M=1.0 
C699 65 86  221.5944E-18 M=1.0 
C700 65 76  55.93725E-18 M=1.0 
C701 65 72  345.2904E-18 M=1.0 
C702 65 70  55.93725E-18 M=1.0 
C703 65 66  55.3986E-18 M=1.0 
C704 64 108  201.6873E-18 M=1.0 
C705 64 71  342.873E-18 M=1.0 
C706 28 84  110.7972E-18 M=1.0 
C707 28 76  110.7972E-18 M=1.0 
C708 28 70  55.3986000000001E-18 M=1.0 
C709 16 84  110.7972E-18 M=1.0 
C710 16 76  110.7972E-18 M=1.0 
C711 16 70  55.3986E-18 M=1.0 
C712 16 28  110.7972E-18 M=1.0 
C713 9 87  55.3986E-18 M=1.0 
C714 9 65  55.3986E-18 M=1.0 
C715 8 87  55.3986E-18 M=1.0 
C716 8 86  55.3986E-18 M=1.0 
C717 8 84  55.3986E-18 M=1.0 
C718 8 76  55.3986E-18 M=1.0 
C719 8 70  55.3986E-18 M=1.0 
C720 8 66  221.5944E-18 M=1.0 
C721 8 65  55.3986E-18 M=1.0 
C722 8 9  311.0229E-18 M=1.0 
C723 2 84  110.7972E-18 M=1.0 
C724 2 76  110.7972E-18 M=1.0 
C725 2 70  55.3986E-18 M=1.0 
C726 2 28  110.7972E-18 M=1.0 
C727 1 84  110.7972E-18 M=1.0 
C728 1 76  110.7972E-18 M=1.0 
C729 1 70  55.3986E-18 M=1.0 
C730 1 16  110.7972E-18 M=1.0 
C731 1 2  110.7972E-18 M=1.0 
C732 VDD 72  34.9776E-18 M=1.0 
C733 VDD 71  34.9776E-18 M=1.0 
C734 VDD 65  1.0735866E-15 M=1.0 
C735 VDD 64  65.5065E-18 M=1.0 
C736 VDD 15  34.9776E-18 M=1.0 
C737 VDD 14  34.9776E-18 M=1.0 
C738 VDD 8  445.7412E-18 M=1.0 
C739 VDD 7  65.5065E-18 M=1.0 
C740 VDD A1  55.3986000000001E-18 M=1.0 
C741 GND 93  4.7994795E-15 M=1.0 
C742 GND 84  4.247406E-15 M=1.0 
C743 GND 72  57.4344E-18 M=1.0 
C744 GND 71  49.167E-18 M=1.0 
C745 GND 65  1.0176642E-15 M=1.0 
C746 GND 64  222.9867E-18 M=1.0 
C747 GND 8  2.6106372E-15 M=1.0 
C748 GND VDD  32.52697155E-15 M=1.0 
C749 CLK 71  90.3762E-18 M=1.0 
C750 CLK 64  143.21295E-18 M=1.0 
C751 CLK VDD  1.32828435E-15 M=1.0 
C752 84 110  209.2176E-18 M=1.0 
C753 76 110  104.6088E-18 M=1.0 
C754 70 110  104.6088E-18 M=1.0 
C755 64 108  69.4476E-18 M=1.0 
C756 28 110  104.6088E-18 M=1.0 
C757 16 110  104.6088E-18 M=1.0 
C758 2 110  104.6088E-18 M=1.0 
C759 GND 110  2.410597575E-15 M=1.0 
C760 GND 108  1.128732075E-15 M=1.0 
C761 CLK 71  52.3044000000001E-18 M=1.0 
C762 CLK 64  94.4298E-18 M=1.0 
C763 VDD 86  129.6405E-18 M=1.0 
C764 VDD 9  62.8560000000001E-18 M=1.0 
C765 GND 87  204.282E-18 M=1.0 
C766 GND 66  166.5684E-18 M=1.0 
C767 GND 65  350.422200000001E-18 M=1.0 
C768 GND 9  147.7116E-18 M=1.0 
C769 28 86  62.3646E-18 M=1.0 
C770 16 87  124.7292E-18 M=1.0 
C771 9 28  124.7292E-18 M=1.0 
C772 9 16  62.3646E-18 M=1.0 
C773 2 66  124.7292E-18 M=1.0 
C774 2 9  62.3646E-18 M=1.0 
C775 1 87  124.7292E-18 M=1.0 
C776 1 66  62.3646E-18 M=1.0 
C777 VDD 86  35.2638E-18 M=1.0 
C778 VDD 65  81.0251999999999E-18 M=1.0 
C779 VDD 28  76.0680000000001E-18 M=1.0 
C780 VDD 16  76.0680000000001E-18 M=1.0 
C781 VDD 9  35.2638E-18 M=1.0 
C782 VDD 2  76.0680000000001E-18 M=1.0 
C783 VDD 1  76.0680000000001E-18 M=1.0 
C784 GND 86  1.0601919E-15 M=1.0 
C785 GND 28  564.3918E-18 M=1.0 
C786 GND 2  757.578599999999E-18 M=1.0 
C787 28 93  110.7972E-18 M=1.0 
C788 28 86  55.93725E-18 M=1.0 
C789 28 66  180.7992E-18 M=1.0 
C790 16 93  110.7972E-18 M=1.0 
C791 16 66  219.384E-18 M=1.0 
C792 9 86  55.3986E-18 M=1.0 
C793 9 66  166.1958E-18 M=1.0 
C794 9 28  55.3986E-18 M=1.0 
C795 9 16  111.33585E-18 M=1.0 
C796 2 93  110.7972E-18 M=1.0 
C797 2 66  55.3986E-18 M=1.0 
C798 2 16  110.7972E-18 M=1.0 
C799 2 9  55.3986E-18 M=1.0 
C800 1 93  110.7972E-18 M=1.0 
C801 1 66  55.3986E-18 M=1.0 
C802 1 28  110.7972E-18 M=1.0 
C803 1 9  55.3986E-18 M=1.0 
C804 VDD 93  1.3095432E-15 M=1.0 
C805 VDD 87  1.3209156E-15 M=1.0 
C806 VDD 86  1.0597788E-15 M=1.0 
C807 VDD 9  204.72975E-18 M=1.0 
C808 VDD 1  1.02615435E-15 M=1.0 
C809 GND 87  669.15E-18 M=1.0 
C810 GND 16  3.21899985E-15 M=1.0 
C811 GND 9  1.666413E-15 M=1.0 
C812 1 110  104.6088E-18 M=1.0 
C813 VDD 7  53.4276000000002E-18 M=1.0 
C814 GND 15  29.8566000000003E-18 M=1.0 
C815 GND 14  29.8566000000001E-18 M=1.0 
C816 GND 8  350.422200000001E-18 M=1.0 
C817 GND 7  182.2824E-18 M=1.0 
C818 15 108  62.3646E-18 M=1.0 
C819 14 108  62.3646000000001E-18 M=1.0 
C820 VDD 108  110.7324E-18 M=1.0 
C821 VDD 15  46.674E-18 M=1.0 
C822 VDD 14  46.6740000000001E-18 M=1.0 
C823 VDD 7  54.2808000000002E-18 M=1.0 
C824 VDD A2  27.1404000000001E-18 M=1.0 
C825 GND 108  219.1122E-18 M=1.0 
C826 GND 15  205.6968E-18 M=1.0 
C827 GND 14  188.6859E-18 M=1.0 
C828 GND 8  707.1354E-18 M=1.0 
C829 GND 7  167.6628E-18 M=1.0 
C830 GND A2  74.6828999999998E-18 M=1.0 
C831 CLK 14  62.3646000000001E-18 M=1.0 
C832 CLK 7  62.3646E-18 M=1.0 
C833 15 108  55.3986E-18 M=1.0 
C834 14 108  75.29535E-18 M=1.0 
C835 8 15  345.2904E-18 M=1.0 
C836 7 108  201.6873E-18 M=1.0 
C837 7 14  342.873E-18 M=1.0 
C838 VDD A2  135.8802E-18 M=1.0 
C839 GND 15  57.4344E-18 M=1.0 
C840 GND 14  49.167E-18 M=1.0 
C841 GND 7  222.9867E-18 M=1.0 
C842 CLK 14  90.3762E-18 M=1.0 
C843 CLK 7  143.21295E-18 M=1.0 
C844 7 108  69.4476E-18 M=1.0 
C845 CLK 108  181.521E-18 M=1.0 
C846 CLK VDD  1.70850465E-15 M=1.0 
C847 VDD 101  26.7138000000002E-18 M=1.0 
C848 GND 101  109.998E-18 M=1.0 
C849 GND 94  39.285E-18 M=1.0 
C850 112 113  62.3646E-18 M=1.0 
C851 101 111  62.3646E-18 M=1.0 
C852 94 112  62.3646E-18 M=1.0 
C853 94 111  62.3646E-18 M=1.0 
C854 87 93  124.7292E-18 M=1.0 
C855 66 93  62.3646E-18 M=1.0 
C856 VDD 113  56.6991E-18 M=1.0 
C857 VDD 112  152.0253E-18 M=1.0 
C858 VDD 101  54.2808E-18 M=1.0 
C859 VDD 94  56.6991E-18 M=1.0 
C860 VDD 93  76.0680000000001E-18 M=1.0 
C861 VDD 3  98.9541E-18 M=1.0 
C862 GND 113  209.3463E-18 M=1.0 
C863 GND 101  176.4513E-18 M=1.0 
C864 GND 94  195.0066E-18 M=1.0 
C865 112 113  55.3986E-18 M=1.0 
C866 101 112  78.3504E-18 M=1.0 
C867 101 111  104.8338E-18 M=1.0 
C868 94 112  50.39325E-18 M=1.0 
C869 94 111  119.3148E-18 M=1.0 
C870 94 101  297.5607E-18 M=1.0 
C871 3 93  233.8533E-18 M=1.0 
C872 VDD 111  2.64360465E-15 M=1.0 
C873 VDD 102  65.5065E-18 M=1.0 
C874 VDD 101  65.5065E-18 M=1.0 
C875 VDD 95  34.9776E-18 M=1.0 
C876 VDD 94  34.9776E-18 M=1.0 
C877 VDD 66  330.2289E-18 M=1.0 
C878 VDD 3  68.5579500000001E-18 M=1.0 
C879 GND 101  157.7223E-18 M=1.0 
C880 GND 94  107.1702E-18 M=1.0 
C881 GND 81  293.6736E-18 M=1.0 
C882 GND 66  1.30877685E-15 M=1.0 
C883 101 112  52.3044E-18 M=1.0 
C884 94 111  37.6677E-18 M=1.0 
C885 93 110  209.2176E-18 M=1.0 
C886 8 110  46.2689999999999E-18 M=1.0 
C887 VDD 110  859.219875E-18 M=1.0 
C888 GND 112  2.35156905E-15 M=1.0 
C889 GND 111  2.07738855E-15 M=1.0 
C890 VDD 108  108.426599999999E-18 M=1.0 
C891 VDD 85  53.4276000000002E-18 M=1.0 
C892 GND 92  29.8566000000003E-18 M=1.0 
C893 GND 91  29.8566000000001E-18 M=1.0 
C894 GND 85  182.2824E-18 M=1.0 
C895 CLK VDD  223.138799999999E-18 M=1.0 
C896 92 108  62.3646E-18 M=1.0 
C897 91 108  62.3646000000001E-18 M=1.0 
C898 VDD 92  46.674E-18 M=1.0 
C899 VDD 91  46.6740000000001E-18 M=1.0 
C900 VDD 85  54.2808000000002E-18 M=1.0 
C901 VDD A0  27.1404000000001E-18 M=1.0 
C902 GND 92  205.6968E-18 M=1.0 
C903 GND 91  188.6859E-18 M=1.0 
C904 GND 85  167.6628E-18 M=1.0 
C905 GND A0  76.5845999999999E-18 M=1.0 
C906 CLK 91  62.3646000000001E-18 M=1.0 
C907 CLK 85  62.3646E-18 M=1.0 
C908 92 108  55.3986E-18 M=1.0 
C909 91 108  75.29535E-18 M=1.0 
C910 86 92  345.2904E-18 M=1.0 
C911 85 108  201.6873E-18 M=1.0 
C912 85 91  342.873E-18 M=1.0 
C913 VDD 108  65.5065E-18 M=1.0 
C914 VDD 92  34.9776E-18 M=1.0 
C915 VDD 91  34.9776E-18 M=1.0 
C916 VDD 85  65.5065E-18 M=1.0 
C917 VDD A0  55.3986000000001E-18 M=1.0 
C918 GND 108  2.77924995E-15 M=1.0 
C919 GND 92  57.4344E-18 M=1.0 
C920 GND 91  49.167E-18 M=1.0 
C921 GND 86  922.5963E-18 M=1.0 
C922 GND 85  222.9867E-18 M=1.0 
C923 CLK 91  90.3762E-18 M=1.0 
C924 CLK 85  143.21295E-18 M=1.0 
C925 CLK GND  81.945E-18 M=1.0 
C926 85 108  69.4476E-18 M=1.0 
C927 VDD 108  1.182449475E-15 M=1.0 
C928 CLK 91  52.3044000000001E-18 M=1.0 
C929 CLK 85  94.4298E-18 M=1.0 
C930 CLK GND  4.4589357E-15 M=1.0 
C931 VDD 162  40.0707E-18 M=1.0 
C932 VDD 152  213.7104E-18 M=1.0 
C933 VDD 146  38.4993E-18 M=1.0 
C934 VDD 145  38.4993E-18 M=1.0 
C935 VDD 144  38.4993E-18 M=1.0 
C936 VDD 142  51.8561999999999E-18 M=1.0 
C937 VDD 141  51.8562000000001E-18 M=1.0 
C938 VDD 140  51.8562E-18 M=1.0 
C939 VDD 134  47.142E-18 M=1.0 
C940 VDD 127  58.1418E-18 M=1.0 
C941 VDD 125  21.2139000000001E-18 M=1.0 
C942 GND 151  222.3531E-18 M=1.0 
C943 GND 146  58.9275E-18 M=1.0 
C944 GND 145  58.9274999999999E-18 M=1.0 
C945 GND 144  58.9275E-18 M=1.0 
C946 GND 142  81.7128000000001E-18 M=1.0 
C947 GND 141  81.7127999999999E-18 M=1.0 
C948 GND 140  81.7128E-18 M=1.0 
C949 150 152  62.3646E-18 M=1.0 
C950 150 151  62.3646E-18 M=1.0 
C951 149 152  62.3646E-18 M=1.0 
C952 149 151  62.3646E-18 M=1.0 
C953 148 152  62.3646E-18 M=1.0 
C954 148 151  62.3646E-18 M=1.0 
C955 147 152  62.3646E-18 M=1.0 
C956 147 151  62.3646E-18 M=1.0 
C957 131 134  62.3646E-18 M=1.0 
C958 129 142  124.7292E-18 M=1.0 
C959 128 131  62.3646E-18 M=1.0 
C960 127 142  62.3646E-18 M=1.0 
C961 125 134  62.3646E-18 M=1.0 
C962 125 131  87.1128E-18 M=1.0 
C963 DFF_OUT_1 134  62.3646E-18 M=1.0 
C964 H_2 145  124.7292E-18 M=1.0 
C965 H_2 141  124.7292E-18 M=1.0 
C966 VDD 162  27.1404E-18 M=1.0 
C967 VDD 158  56.6991E-18 M=1.0 
C968 VDD 152  196.5996E-18 M=1.0 
C969 VDD 146  46.3662E-18 M=1.0 
C970 VDD 145  46.3662E-18 M=1.0 
C971 VDD 144  46.3662E-18 M=1.0 
C972 VDD 142  147.1671E-18 M=1.0 
C973 VDD 138  39.0672E-18 M=1.0 
C974 VDD 128  48.5262E-18 M=1.0 
C975 VDD 122  27.1404E-18 M=1.0 
C976 VDD H_2  99.4158E-18 M=1.0 
C977 VDD OUT_2  47.8611E-18 M=1.0 
C978 H_1 146  124.7292E-18 M=1.0 
C979 H_1 142  124.7292E-18 M=1.0 
C980 H_1 VDD  140.2308E-18 M=1.0 
C981 _DFF_OUT_2 VDD  121.4667E-18 M=1.0 
C982 H_0 144  124.7292E-18 M=1.0 
C983 H_0 140  124.7292E-18 M=1.0 
C984 H_0 VDD  143.8803E-18 M=1.0 
C985 GND 154  119.63115E-18 M=1.0 
C986 GND 150  137.9502E-18 M=1.0 
C987 GND 149  137.9502E-18 M=1.0 
C988 GND 148  137.9502E-18 M=1.0 
C989 GND 147  137.9502E-18 M=1.0 
C990 GND 146  92.3202E-18 M=1.0 
C991 GND 145  92.3202E-18 M=1.0 
C992 GND 144  92.3202E-18 M=1.0 
C993 GND 143  92.3201999999999E-18 M=1.0 
C994 GND 140  151.0308E-18 M=1.0 
C995 GND 139  152.262E-18 M=1.0 
C996 GND 134  448.4826E-18 M=1.0 
C997 GND 131  39.1662E-18 M=1.0 
C998 GND 127  130.167E-18 M=1.0 
C999 GND 125  94.068E-18 M=1.0 
C1000 GND 122  46.1574E-18 M=1.0 
C1001 GND H_2  334.7541E-18 M=1.0 
C1002 GND H_1  268.524E-18 M=1.0 
C1003 GND _DFF_OUT_2  432.1692E-18 M=1.0 
C1004 GND H_0  308.6577E-18 M=1.0 
C1005 DFF_OUT_6 VDD  154.6749E-18 M=1.0 
C1006 DFF_OUT_6 GND  1.1417724E-15 M=1.0 
C1007 DFF_OUT_5 125  105.67395E-18 M=1.0 
C1008 DFF_OUT_5 VDD  75.3093E-18 M=1.0 
C1009 DFF_OUT_5 GND  916.66305E-18 M=1.0 
C1010 DFF_OUT_4 VDD  109.5948E-18 M=1.0 
C1011 DFF_OUT_4 GND  226.34595E-18 M=1.0 
C1012 _DFF_OUT_6 GND  261.2691E-18 M=1.0 
C1013 _DFF_OUT_5 VDD  75.0015E-18 M=1.0 
C1014 _DFF_OUT_5 GND  231.7653E-18 M=1.0 
C1015 DFF_OUT_2 VDD  124.0389E-18 M=1.0 
C1016 DFF_OUT_2 GND  706.8222E-18 M=1.0 
C1017 H_3 143  124.7292E-18 M=1.0 
C1018 H_3 139  124.7292E-18 M=1.0 
C1019 H_3 VDD  137.69145E-18 M=1.0 
C1020 H_3 GND  494.63955E-18 M=1.0 
C1021 152 154  55.3986E-18 M=1.0 
C1022 148 152  34.9776E-18 M=1.0 
C1023 142 146  59.62635E-18 M=1.0 
C1024 141 145  59.62635E-18 M=1.0 
C1025 140 144  59.62635E-18 M=1.0 
C1026 139 143  59.62635E-18 M=1.0 
C1027 128 138  74.691E-18 M=1.0 
C1028 128 134  90.3762E-18 M=1.0 
C1029 128 131  100.4841E-18 M=1.0 
C1030 125 131  34.9776E-18 M=1.0 
C1031 125 128  120.9051E-18 M=1.0 
C1032 122 125  55.3986E-18 M=1.0 
C1033 _DFF_OUT_4 146  145.0206E-18 M=1.0 
C1034 _DFF_OUT_4 142  250.29945E-18 M=1.0 
C1035 _DFF_OUT_4 138  110.1303E-18 M=1.0 
C1036 _DFF_OUT_4 129  34.9776E-18 M=1.0 
C1037 _DFF_OUT_4 128  34.9776E-18 M=1.0 
C1038 _DFF_OUT_4 127  34.9776E-18 M=1.0 
C1039 H_2 145  55.3986E-18 M=1.0 
C1040 H_2 141  65.42955E-18 M=1.0 
C1041 VDD 146  250.4286E-18 M=1.0 
C1042 VDD 145  250.4286E-18 M=1.0 
C1043 VDD 144  250.4286E-18 M=1.0 
C1044 VDD 143  250.4286E-18 M=1.0 
C1045 VDD 128  488.2302E-18 M=1.0 
C1046 VDD 127  797.38335E-18 M=1.0 
C1047 VDD 125  130.5198E-18 M=1.0 
C1048 VDD H_2  135.8802E-18 M=1.0 
C1049 H_1 146  55.3986E-18 M=1.0 
C1050 H_1 142  65.42955E-18 M=1.0 
C1051 H_1 VDD  135.8802E-18 M=1.0 
C1052 _DFF_OUT_2 144  55.3986E-18 M=1.0 
C1053 _DFF_OUT_2 140  65.42955E-18 M=1.0 
C1054 H_0 144  55.3986E-18 M=1.0 
C1055 H_0 140  65.42955E-18 M=1.0 
C1056 H_0 VDD  104.5971E-18 M=1.0 
C1057 GND 165  137.0394E-18 M=1.0 
C1058 GND 146  252.9216E-18 M=1.0 
C1059 GND 145  252.9216E-18 M=1.0 
C1060 GND 144  252.9216E-18 M=1.0 
C1061 GND 143  252.9216E-18 M=1.0 
C1062 GND 142  346.2345E-18 M=1.0 
C1063 GND 141  346.2345E-18 M=1.0 
C1064 GND 140  346.2345E-18 M=1.0 
C1065 GND 139  346.2345E-18 M=1.0 
C1066 GND 128  852.8643E-18 M=1.0 
C1067 GND 125  74.1006E-18 M=1.0 
C1068 DFF_OUT_6 GND  1.4821425E-15 M=1.0 
C1069 DFF_OUT_5 134  125.3538E-18 M=1.0 
C1070 DFF_OUT_5 131  100.4841E-18 M=1.0 
C1071 DFF_OUT_5 128  65.9682E-18 M=1.0 
C1072 DFF_OUT_5 125  119.3634E-18 M=1.0 
C1073 DFF_OUT_5 122  65.9682E-18 M=1.0 
C1074 DFF_OUT_5 VDD  451.7415E-18 M=1.0 
C1075 DFF_OUT_5 GND  1.9103049E-15 M=1.0 
C1076 DFF_OUT_4 VDD  210.2778E-18 M=1.0 
C1077 DFF_OUT_4 GND  3.8796444E-15 M=1.0 
C1078 _DFF_OUT_6 143  55.3986E-18 M=1.0 
C1079 _DFF_OUT_6 139  65.42955E-18 M=1.0 
C1080 _DFF_OUT_5 145  55.3986E-18 M=1.0 
C1081 _DFF_OUT_5 141  65.42955E-18 M=1.0 
C1082 _DFF_OUT_5 VDD  1.5475599E-15 M=1.0 
C1083 _DFF_OUT_5 GND  3.4379973E-15 M=1.0 
C1084 DFF_OUT_2 GND  2.214288E-15 M=1.0 
C1085 H_3 143  55.3986E-18 M=1.0 
C1086 H_3 139  65.42955E-18 M=1.0 
C1087 H_3 VDD  135.8802E-18 M=1.0 
C1088 151 152  706.2894E-18 M=1.0 
C1089 150 152  37.6677E-18 M=1.0 
C1090 149 152  37.6677E-18 M=1.0 
C1091 148 152  37.6677E-18 M=1.0 
C1092 147 152  37.6677E-18 M=1.0 
C1093 142 146  130.1292E-18 M=1.0 
C1094 141 145  130.1292E-18 M=1.0 
C1095 140 144  130.1292E-18 M=1.0 
C1096 139 143  130.1292E-18 M=1.0 
C1097 129 142  37.6677E-18 M=1.0 
C1098 129 140  37.6677E-18 M=1.0 
C1099 128 138  114.8985E-18 M=1.0 
C1100 127 142  75.1248E-18 M=1.0 
C1101 127 128  189.8829E-18 M=1.0 
C1102 _DFF_OUT_4 129  52.3044E-18 M=1.0 
C1103 _DFF_OUT_4 128  104.6088E-18 M=1.0 
C1104 _DFF_OUT_4 127  52.3044E-18 M=1.0 
C1105 H_2 145  37.6677E-18 M=1.0 
C1106 VDD 152  1.1372994E-15 M=1.0 
C1107 VDD 151  493.8219E-18 M=1.0 
C1108 VDD 146  52.3044E-18 M=1.0 
C1109 VDD 145  52.3044E-18 M=1.0 
C1110 VDD 144  52.3044E-18 M=1.0 
C1111 VDD 143  52.3044E-18 M=1.0 
C1112 VDD 142  52.3044E-18 M=1.0 
C1113 VDD 141  52.3044E-18 M=1.0 
C1114 VDD 140  52.3044E-18 M=1.0 
C1115 VDD 139  52.3044E-18 M=1.0 
C1116 VDD 129  640.033875E-18 M=1.0 
C1117 VDD 128  235.9845E-18 M=1.0 
C1118 H_1 146  37.6677E-18 M=1.0 
C1119 _DFF_OUT_2 129  52.3044E-18 M=1.0 
C1120 _DFF_OUT_2 128  104.6088E-18 M=1.0 
C1121 H_0 144  37.6677E-18 M=1.0 
C1122 GND 152  2.99562525E-15 M=1.0 
C1123 GND 146  278.2449E-18 M=1.0 
C1124 GND 145  278.2449E-18 M=1.0 
C1125 GND 144  278.2449E-18 M=1.0 
C1126 GND 143  278.2449E-18 M=1.0 
C1127 GND VDD  4.7622015E-15 M=1.0 
C1128 DFF_OUT_6 125  52.3044E-18 M=1.0 
C1129 DFF_OUT_6 122  155.8368E-18 M=1.0 
C1130 DFF_OUT_6 VDD  526.8573E-18 M=1.0 
C1131 DFF_OUT_5 134  33.6204E-18 M=1.0 
C1132 DFF_OUT_5 129  52.3044E-18 M=1.0 
C1133 DFF_OUT_5 128  104.6088E-18 M=1.0 
C1134 DFF_OUT_5 127  52.3044E-18 M=1.0 
C1135 DFF_OUT_5 _DFF_OUT_4  104.6088E-18 M=1.0 
C1136 DFF_OUT_5 VDD  218.925675E-18 M=1.0 
C1137 DFF_OUT_5 _DFF_OUT_2  52.3044E-18 M=1.0 
C1138 DFF_OUT_5 DFF_OUT_6  52.3044E-18 M=1.0 
C1139 DFF_OUT_4 129  52.3044E-18 M=1.0 
C1140 DFF_OUT_4 DFF_OUT_5  52.3044E-18 M=1.0 
C1141 _DFF_OUT_6 128  187.6248E-18 M=1.0 
C1142 _DFF_OUT_6 DFF_OUT_5  164.53305E-18 M=1.0 
C1143 _DFF_OUT_5 125  70.614E-18 M=1.0 
C1144 _DFF_OUT_5 DFF_OUT_5  52.3044E-18 M=1.0 
C1145 DFF_OUT_2 144  173.0178E-18 M=1.0 
C1146 DFF_OUT_2 142  159.57315E-18 M=1.0 
C1147 DFF_OUT_2 140  52.3044E-18 M=1.0 
C1148 DFF_OUT_2 129  52.3044E-18 M=1.0 
C1149 DFF_OUT_2 _DFF_OUT_4  52.3044E-18 M=1.0 
C1150 DFF_OUT_2 VDD  577.69785E-18 M=1.0 
C1151 DFF_OUT_2 _DFF_OUT_2  104.6088E-18 M=1.0 
C1152 DFF_OUT_2 GND  1.27809585E-15 M=1.0 
C1153 DFF_OUT_2 DFF_OUT_5  52.3044E-18 M=1.0 
C1154 H_3 143  37.6677E-18 M=1.0 
C1155 VDD 135  47.142E-18 M=1.0 
C1156 VDD 129  58.1418E-18 M=1.0 
C1157 VDD 126  21.2139E-18 M=1.0 
C1158 _DFF_OUT_3 VDD  53.4276E-18 M=1.0 
C1159 GND 138  43.2135E-18 M=1.0 
C1160 GND 136  43.2135E-18 M=1.0 
C1161 GND 135  66.7845E-18 M=1.0 
C1162 GND 134  66.7845E-18 M=1.0 
C1163 GND 132  58.9275E-18 M=1.0 
C1164 GND 131  58.9275000000001E-18 M=1.0 
C1165 GND 129  174.4254E-18 M=1.0 
C1166 GND 127  127.2834E-18 M=1.0 
C1167 GND 126  27.4995E-18 M=1.0 
C1168 GND 125  27.4995E-18 M=1.0 
C1169 DFF_OUT_5 VDD  155.96145E-18 M=1.0 
C1170 DFF_OUT_5 GND  73.46295E-18 M=1.0 
C1171 DFF_OUT_3 VDD  65.2131E-18 M=1.0 
C1172 DFF_OUT_3 GND  52.6419E-18 M=1.0 
C1173 _DFF_OUT_5 VDD  77.7843000000001E-18 M=1.0 
C1174 _DFF_OUT_5 GND  252.9954E-18 M=1.0 
C1175 132 135  62.3646E-18 M=1.0 
C1176 129 132  62.3646E-18 M=1.0 
C1177 128 140  124.7292E-18 M=1.0 
C1178 127 140  62.3646E-18 M=1.0 
C1179 126 135  62.3646E-18 M=1.0 
C1180 126 132  87.1128E-18 M=1.0 
C1181 VDD 140  147.1671E-18 M=1.0 
C1182 VDD 136  39.0672E-18 M=1.0 
C1183 VDD 135  69.4944E-18 M=1.0 
C1184 VDD 129  38.99025E-18 M=1.0 
C1185 VDD 126  151.3224E-18 M=1.0 
C1186 VDD 123  27.1404E-18 M=1.0 
C1187 _DFF_OUT_3 135  62.3646E-18 M=1.0 
C1188 GND 142  151.0308E-18 M=1.0 
C1189 GND 138  75.6612E-18 M=1.0 
C1190 GND 136  156.58695E-18 M=1.0 
C1191 GND 135  448.4826E-18 M=1.0 
C1192 GND 132  39.1662E-18 M=1.0 
C1193 GND 126  94.068E-18 M=1.0 
C1194 GND 123  46.1574E-18 M=1.0 
C1195 GND _DFF_OUT_4  267.0786E-18 M=1.0 
C1196 GND _DFF_OUT_3  525.5946E-18 M=1.0 
C1197 DFF_OUT_5 126  105.67395E-18 M=1.0 
C1198 DFF_OUT_4 _DFF_OUT_3  62.3646E-18 M=1.0 
C1199 DFF_OUT_3 135  62.3646E-18 M=1.0 
C1200 DFF_OUT_3 _DFF_OUT_4  62.3646E-18 M=1.0 
C1201 DFF_OUT_3 VDD  32.6421E-18 M=1.0 
C1202 DFF_OUT_3 GND  371.5074E-18 M=1.0 
C1203 _DFF_OUT_5 126  62.3646E-18 M=1.0 
C1204 _DFF_OUT_5 DFF_OUT_6  124.7292E-18 M=1.0 
C1205 129 136  20.7792E-18 M=1.0 
C1206 129 135  90.3762E-18 M=1.0 
C1207 129 132  100.40715E-18 M=1.0 
C1208 128 140  166.1958E-18 M=1.0 
C1209 128 136  34.9776E-18 M=1.0 
C1210 128 129  20.7792E-18 M=1.0 
C1211 127 129  20.7792E-18 M=1.0 
C1212 127 128  34.9776E-18 M=1.0 
C1213 126 132  34.9776E-18 M=1.0 
C1214 126 129  120.82815E-18 M=1.0 
C1215 123 126  55.3986E-18 M=1.0 
C1216 _DFF_OUT_4 134  113.2758E-18 M=1.0 
C1217 VDD 126  130.5198E-18 M=1.0 
C1218 VDD _DFF_OUT_4  1.2171519E-15 M=1.0 
C1219 _DFF_OUT_3 _DFF_OUT_4  55.3986E-18 M=1.0 
C1220 GND 129  1.2261537E-15 M=1.0 
C1221 GND 126  74.1006E-18 M=1.0 
C1222 GND _DFF_OUT_4  2.7010089E-15 M=1.0 
C1223 DFF_OUT_5 _DFF_OUT_4  55.3986E-18 M=1.0 
C1224 DFF_OUT_5 _DFF_OUT_3  55.3986E-18 M=1.0 
C1225 DFF_OUT_4 142  60.46875E-18 M=1.0 
C1226 DFF_OUT_4 138  34.9776E-18 M=1.0 
C1227 DFF_OUT_4 135  60.165E-18 M=1.0 
C1228 DFF_OUT_4 129  34.9776E-18 M=1.0 
C1229 DFF_OUT_4 127  34.9776E-18 M=1.0 
C1230 _DFF_OUT_6 126  89.48835E-18 M=1.0 
C1231 _DFF_OUT_6 DFF_OUT_6  171.26595E-18 M=1.0 
C1232 _DFF_OUT_6 DFF_OUT_5  133.3746E-18 M=1.0 
C1233 DFF_OUT_3 135  55.3986E-18 M=1.0 
C1234 DFF_OUT_3 134  299.3148E-18 M=1.0 
C1235 DFF_OUT_3 _DFF_OUT_3  187.5924E-18 M=1.0 
C1236 DFF_OUT_3 GND  1.0568331E-15 M=1.0 
C1237 DFF_OUT_3 DFF_OUT_5  55.3986E-18 M=1.0 
C1238 DFF_OUT_3 DFF_OUT_4  258.642E-18 M=1.0 
C1239 _DFF_OUT_5 DFF_OUT_6  131.2866E-18 M=1.0 
C1240 127 140  75.6513E-18 M=1.0 
C1241 VDD 127  219.86595E-18 M=1.0 
C1242 VDD _DFF_OUT_4  189.830025E-18 M=1.0 
C1243 _DFF_OUT_3 VDD  52.3044E-18 M=1.0 
C1244 _DFF_OUT_2 _DFF_OUT_4  52.3044E-18 M=1.0 
C1245 GND 140  44.1036E-18 M=1.0 
C1246 GND 138  37.6677E-18 M=1.0 
C1247 GND 136  192.4263E-18 M=1.0 
C1248 GND 127  1.218818925E-15 M=1.0 
C1249 GND _DFF_OUT_4  2.242333575E-15 M=1.0 
C1250 DFF_OUT_6 _DFF_OUT_3  52.3044E-18 M=1.0 
C1251 DFF_OUT_6 GND  639.31725E-18 M=1.0 
C1252 DFF_OUT_5 _DFF_OUT_3  52.3044E-18 M=1.0 
C1253 DFF_OUT_5 GND  392.5071E-18 M=1.0 
C1254 DFF_OUT_4 128  153.4293E-18 M=1.0 
C1255 DFF_OUT_4 127  104.6088E-18 M=1.0 
C1256 DFF_OUT_4 _DFF_OUT_4  156.9132E-18 M=1.0 
C1257 DFF_OUT_4 VDD  312.459525E-18 M=1.0 
C1258 DFF_OUT_4 _DFF_OUT_2  156.9132E-18 M=1.0 
C1259 DFF_OUT_4 GND  1.3126095E-15 M=1.0 
C1260 _DFF_OUT_6 126  150.1443E-18 M=1.0 
C1261 _DFF_OUT_6 VDD  368.2359E-18 M=1.0 
C1262 _DFF_OUT_6 _DFF_OUT_3  52.3044E-18 M=1.0 
C1263 DFF_OUT_3 VDD  52.3044E-18 M=1.0 
C1264 DFF_OUT_3 DFF_OUT_6  52.3044E-18 M=1.0 
C1265 DFF_OUT_3 DFF_OUT_5  52.3044E-18 M=1.0 
C1266 DFF_OUT_3 DFF_OUT_4  227.9799E-18 M=1.0 
C1267 DFF_OUT_3 _DFF_OUT_6  52.3044E-18 M=1.0 
C1268 _DFF_OUT_5 _DFF_OUT_4  52.3044E-18 M=1.0 
C1269 _DFF_OUT_5 _DFF_OUT_3  52.3044E-18 M=1.0 
C1270 _DFF_OUT_5 _DFF_OUT_6  140.1714E-18 M=1.0 
C1271 _DFF_OUT_5 DFF_OUT_3  52.3044E-18 M=1.0 
C1272 VDD 133  47.1419999999999E-18 M=1.0 
C1273 VDD 124  21.2139E-18 M=1.0 
C1274 VDD DFF_OUT_1  57.945375E-18 M=1.0 
C1275 DFF_OUT_0 VDD  57.9453750000001E-18 M=1.0 
C1276 _DFF_OUT_1 VDD  53.4276000000001E-18 M=1.0 
C1277 GND 139  81.7127999999999E-18 M=1.0 
C1278 GND 137  43.2135E-18 M=1.0 
C1279 GND 133  66.7845000000001E-18 M=1.0 
C1280 GND 130  58.9275000000004E-18 M=1.0 
C1281 GND 128  136.7118E-18 M=1.0 
C1282 GND 124  27.4995000000001E-18 M=1.0 
C1283 GND DFF_OUT_1  59.9096249999999E-18 M=1.0 
C1284 GND DFF_OUT_0  59.909625E-18 M=1.0 
C1285 GND _DFF_OUT_1  206.6391E-18 M=1.0 
C1286 _DFF_OUT_0 VDD  53.4276000000002E-18 M=1.0 
C1287 DFF_OUT_4 VDD  78.5699999999998E-18 M=1.0 
C1288 130 133  62.3646E-18 M=1.0 
C1289 129 141  124.7292E-18 M=1.0 
C1290 129 139  124.7292E-18 M=1.0 
C1291 128 141  62.3646E-18 M=1.0 
C1292 128 139  62.3646E-18 M=1.0 
C1293 127 130  62.3646E-18 M=1.0 
C1294 124 133  62.3646E-18 M=1.0 
C1295 124 130  87.1128E-18 M=1.0 
C1296 _DFF_OUT_4 124  62.3646E-18 M=1.0 
C1297 VDD 141  147.1671E-18 M=1.0 
C1298 VDD 139  147.5298E-18 M=1.0 
C1299 VDD 137  39.0672E-18 M=1.0 
C1300 VDD 134  69.4944E-18 M=1.0 
C1301 VDD 133  69.4944E-18 M=1.0 
C1302 VDD 127  41.6889E-18 M=1.0 
C1303 VDD 125  151.3224E-18 M=1.0 
C1304 VDD 124  151.3224E-18 M=1.0 
C1305 VDD 121  27.1404E-18 M=1.0 
C1306 VDD _DFF_OUT_4  102.1419E-18 M=1.0 
C1307 DFF_OUT_0 133  62.3646E-18 M=1.0 
C1308 _DFF_OUT_2 DFF_OUT_1  62.3646E-18 M=1.0 
C1309 _DFF_OUT_1 134  62.3646E-18 M=1.0 
C1310 GND 141  151.0308E-18 M=1.0 
C1311 GND 137  75.6612E-18 M=1.0 
C1312 GND 130  39.1662E-18 M=1.0 
C1313 GND 129  185.83875E-18 M=1.0 
C1314 GND 128  156.2247E-18 M=1.0 
C1315 GND 121  46.1574E-18 M=1.0 
C1316 GND _DFF_OUT_1  170.2845E-18 M=1.0 
C1317 _DFF_OUT_0 133  62.3646E-18 M=1.0 
C1318 DFF_OUT_6 _DFF_OUT_4  62.3646E-18 M=1.0 
C1319 DFF_OUT_4 124  105.67395E-18 M=1.0 
C1320 _DFF_OUT_6 DFF_OUT_5  304.884E-18 M=1.0 
C1321 _DFF_OUT_5 125  62.3646E-18 M=1.0 
C1322 DFF_OUT_2 _DFF_OUT_1  62.3646E-18 M=1.0 
C1323 128 137  114.4917E-18 M=1.0 
C1324 127 133  90.3762E-18 M=1.0 
C1325 127 130  100.40715E-18 M=1.0 
C1326 124 130  34.9776E-18 M=1.0 
C1327 124 127  120.82815E-18 M=1.0 
C1328 121 124  55.3986E-18 M=1.0 
C1329 DFF_OUT_1 134  73.8648E-18 M=1.0 
C1330 VDD 133  55.3986E-18 M=1.0 
C1331 VDD 124  130.5198E-18 M=1.0 
C1332 VDD DFF_OUT_1  47.74545E-18 M=1.0 
C1333 _DFF_OUT_2 DFF_OUT_1  55.3986E-18 M=1.0 
C1334 GND 127  576.7623E-18 M=1.0 
C1335 GND 124  74.1006E-18 M=1.0 
C1336 GND DFF_OUT_1  43.10865E-18 M=1.0 
C1337 _DFF_OUT_0 124  133.87995E-18 M=1.0 
C1338 _DFF_OUT_0 _DFF_OUT_4  59.436E-18 M=1.0 
C1339 _DFF_OUT_0 VDD  192.4776E-18 M=1.0 
C1340 DFF_OUT_6 133  125.3538E-18 M=1.0 
C1341 DFF_OUT_6 130  100.4841E-18 M=1.0 
C1342 DFF_OUT_6 127  65.9682E-18 M=1.0 
C1343 DFF_OUT_6 124  65.5065E-18 M=1.0 
C1344 DFF_OUT_6 121  85.6575E-18 M=1.0 
C1345 DFF_OUT_6 VDD  245.3391E-18 M=1.0 
C1346 DFF_OUT_6 _DFF_OUT_0  134.75475E-18 M=1.0 
C1347 DFF_OUT_4 133  380.68425E-18 M=1.0 
C1348 _DFF_OUT_6 125  65.2635E-18 M=1.0 
C1349 _DFF_OUT_6 124  65.2635E-18 M=1.0 
C1350 _DFF_OUT_6 _DFF_OUT_4  49.176E-18 M=1.0 
C1351 _DFF_OUT_6 DFF_OUT_4  49.1985E-18 M=1.0 
C1352 _DFF_OUT_5 137  75.1527E-18 M=1.0 
C1353 _DFF_OUT_5 127  34.9776E-18 M=1.0 
C1354 _DFF_OUT_5 _DFF_OUT_6  98.352E-18 M=1.0 
C1355 DFF_OUT_2 134  94.2021E-18 M=1.0 
C1356 DFF_OUT_2 133  60.165E-18 M=1.0 
C1357 DFF_OUT_2 DFF_OUT_1  144.1728E-18 M=1.0 
C1358 DFF_OUT_2 VDD  251.1774E-18 M=1.0 
C1359 DFF_OUT_2 DFF_OUT_0  49.176E-18 M=1.0 
C1360 129 141  148.71645E-18 M=1.0 
C1361 129 137  51.0561E-18 M=1.0 
C1362 128 137  111.78585E-18 M=1.0 
C1363 128 129  25.6374E-18 M=1.0 
C1364 _DFF_OUT_2 127  104.6088E-18 M=1.0 
C1365 _DFF_OUT_2 DFF_OUT_1  194.900625E-18 M=1.0 
C1366 _DFF_OUT_2 VDD  122.9121E-18 M=1.0 
C1367 _DFF_OUT_1 133  93.7305E-18 M=1.0 
C1368 _DFF_OUT_1 130  141.3855E-18 M=1.0 
C1369 _DFF_OUT_1 127  52.3044E-18 M=1.0 
C1370 _DFF_OUT_1 VDD  307.445175E-18 M=1.0 
C1371 GND 137  37.6677E-18 M=1.0 
C1372 GND 129  1.780714575E-15 M=1.0 
C1373 GND 128  1.1781747E-15 M=1.0 
C1374 GND _DFF_OUT_2  1.52013015E-15 M=1.0 
C1375 GND _DFF_OUT_1  1.272761775E-15 M=1.0 
C1376 _DFF_OUT_0 _DFF_OUT_4  52.3044E-18 M=1.0 
C1377 DFF_OUT_6 129  52.3044E-18 M=1.0 
C1378 DFF_OUT_6 128  52.3044E-18 M=1.0 
C1379 DFF_OUT_6 127  52.3044E-18 M=1.0 
C1380 DFF_OUT_6 124  52.3044E-18 M=1.0 
C1381 DFF_OUT_6 121  141.435E-18 M=1.0 
C1382 DFF_OUT_6 _DFF_OUT_4  57.4173E-18 M=1.0 
C1383 DFF_OUT_6 _DFF_OUT_2  52.3044E-18 M=1.0 
C1384 DFF_OUT_6 _DFF_OUT_1  52.3044E-18 M=1.0 
C1385 DFF_OUT_6 _DFF_OUT_0  119.8719E-18 M=1.0 
C1386 DFF_OUT_5 125  211.584825E-18 M=1.0 
C1387 DFF_OUT_4 124  231.738075E-18 M=1.0 
C1388 DFF_OUT_4 DFF_OUT_1  51.138E-18 M=1.0 
C1389 DFF_OUT_4 _DFF_OUT_1  52.3044E-18 M=1.0 
C1390 DFF_OUT_4 DFF_OUT_6  104.6088E-18 M=1.0 
C1391 _DFF_OUT_6 127  187.6248E-18 M=1.0 
C1392 _DFF_OUT_6 125  252.9882E-18 M=1.0 
C1393 _DFF_OUT_6 124  181.39725E-18 M=1.0 
C1394 _DFF_OUT_6 _DFF_OUT_4  86.9805E-18 M=1.0 
C1395 _DFF_OUT_6 GND  694.307475E-18 M=1.0 
C1396 _DFF_OUT_6 _DFF_OUT_0  128.8809E-18 M=1.0 
C1397 _DFF_OUT_6 DFF_OUT_6  52.3044E-18 M=1.0 
C1398 _DFF_OUT_6 DFF_OUT_4  136.78245E-18 M=1.0 
C1399 _DFF_OUT_5 129  52.3044E-18 M=1.0 
C1400 _DFF_OUT_5 128  132.0732E-18 M=1.0 
C1401 _DFF_OUT_5 127  52.3044E-18 M=1.0 
C1402 _DFF_OUT_5 VDD  530.63775E-18 M=1.0 
C1403 _DFF_OUT_5 _DFF_OUT_2  52.3044E-18 M=1.0 
C1404 _DFF_OUT_5 _DFF_OUT_1  52.3044E-18 M=1.0 
C1405 _DFF_OUT_5 GND  817.0281E-18 M=1.0 
C1406 _DFF_OUT_5 DFF_OUT_6  114.8346E-18 M=1.0 
C1407 _DFF_OUT_5 DFF_OUT_4  52.3044E-18 M=1.0 
C1408 DFF_OUT_2 133  56.3436E-18 M=1.0 
C1409 DFF_OUT_2 128  52.3044E-18 M=1.0 
C1410 DFF_OUT_2 127  104.6088E-18 M=1.0 
C1411 DFF_OUT_2 DFF_OUT_0  51.110775E-18 M=1.0 
C1412 DFF_OUT_2 _DFF_OUT_1  180.868725E-18 M=1.0 
C1413 DFF_OUT_2 DFF_OUT_6  52.3044E-18 M=1.0 
C1414 DFF_OUT_2 DFF_OUT_4  156.9132E-18 M=1.0 
C1415 DFF_OUT_2 _DFF_OUT_5  52.3044E-18 M=1.0 
C1416 DFF_OUT_1 134  87.12585E-18 M=1.0 
C1417 DFF_OUT_1 127  49.5477E-18 M=1.0 
C1418 VDD DFF_OUT_1  179.4771E-18 M=1.0 
C1419 GND DFF_OUT_1  823.8654E-18 M=1.0 
C1420 _DFF_OUT_0 DFF_OUT_1  75.5973E-18 M=1.0 
C1421 DFF_OUT_6 DFF_OUT_1  49.5477E-18 M=1.0 
C1422 DFF_OUT_4 DFF_OUT_1  49.5477E-18 M=1.0 
C1423 _DFF_OUT_5 DFF_OUT_1  49.5477E-18 M=1.0 
C1424 VDD 164  40.0707E-18 M=1.0 
C1425 VDD 163  40.0707E-18 M=1.0 
C1426 VDD 151  146.9259E-18 M=1.0 
C1427 GND 164  148.4973E-18 M=1.0 
C1428 GND 163  148.4973E-18 M=1.0 
C1429 GND 160  38.4993E-18 M=1.0 
C1430 GND 159  38.4993E-18 M=1.0 
C1431 GND 152  128.8548E-18 M=1.0 
C1432 GND 150  38.4993E-18 M=1.0 
C1433 GND 149  38.4993E-18 M=1.0 
C1434 152 156  62.3646E-18 M=1.0 
C1435 152 155  62.3646E-18 M=1.0 
C1436 151 160  62.3646E-18 M=1.0 
C1437 151 159  62.3646E-18 M=1.0 
C1438 VDD 164  27.1404E-18 M=1.0 
C1439 VDD 163  27.1404E-18 M=1.0 
C1440 VDD 160  56.6991E-18 M=1.0 
C1441 VDD 159  56.6991E-18 M=1.0 
C1442 VDD 156  54.2808E-18 M=1.0 
C1443 VDD 155  54.2808E-18 M=1.0 
C1444 VDD 151  67.0428E-18 M=1.0 
C1445 OUT_1 VDD  47.8611E-18 M=1.0 
C1446 OUT_0 VDD  47.8611E-18 M=1.0 
C1447 GND 164  162.0072E-18 M=1.0 
C1448 GND 163  162.0072E-18 M=1.0 
C1449 GND 160  226.4616E-18 M=1.0 
C1450 GND 159  226.4616E-18 M=1.0 
C1451 GND 156  119.63115E-18 M=1.0 
C1452 GND 155  119.63115E-18 M=1.0 
C1453 GND OUT_1  98.3826E-18 M=1.0 
C1454 GND OUT_0  98.3826E-18 M=1.0 
C1455 160 164  306.8514E-18 M=1.0 
C1456 159 163  306.8514E-18 M=1.0 
C1457 152 156  55.3986E-18 M=1.0 
C1458 152 155  55.3986E-18 M=1.0 
C1459 151 160  120.9051E-18 M=1.0 
C1460 151 159  120.9051E-18 M=1.0 
C1461 151 156  224.6967E-18 M=1.0 
C1462 151 155  224.6967E-18 M=1.0 
C1463 151 152  139.9104E-18 M=1.0 
C1464 150 152  34.9776E-18 M=1.0 
C1465 150 151  65.31255E-18 M=1.0 
C1466 149 152  34.9776E-18 M=1.0 
C1467 149 151  65.31255E-18 M=1.0 
C1468 OUT_1 163  55.3986E-18 M=1.0 
C1469 OUT_0 164  55.3986E-18 M=1.0 
C1470 GND 164  559.068525E-18 M=1.0 
C1471 GND 163  559.068525E-18 M=1.0 
C1472 GND 160  113.0463E-18 M=1.0 
C1473 GND 159  113.0463E-18 M=1.0 
C1474 150 151  223.1748E-18 M=1.0 
C1475 149 151  223.1748E-18 M=1.0 
C1476 VDD 161  40.0707E-18 M=1.0 
C1477 GND 162  148.4973E-18 M=1.0 
C1478 GND 161  148.4973E-18 M=1.0 
C1479 GND 158  38.4993E-18 M=1.0 
C1480 GND 157  38.4993000000001E-18 M=1.0 
C1481 GND 148  38.4993E-18 M=1.0 
C1482 GND 147  38.4993E-18 M=1.0 
C1483 152 154  62.3646E-18 M=1.0 
C1484 152 153  62.3646E-18 M=1.0 
C1485 151 158  62.3646E-18 M=1.0 
C1486 151 157  62.3646E-18 M=1.0 
C1487 VDD 161  27.1404E-18 M=1.0 
C1488 VDD 157  56.6991E-18 M=1.0 
C1489 VDD 154  54.2808E-18 M=1.0 
C1490 VDD 153  54.2808E-18 M=1.0 
C1491 GND 162  162.0072E-18 M=1.0 
C1492 GND 161  162.0072E-18 M=1.0 
C1493 GND 158  226.4616E-18 M=1.0 
C1494 GND 157  226.4616E-18 M=1.0 
C1495 GND 153  119.63115E-18 M=1.0 
C1496 GND 151  339.9138E-18 M=1.0 
C1497 GND OUT_2  98.3826E-18 M=1.0 
C1498 OUT_3 VDD  47.8611E-18 M=1.0 
C1499 OUT_3 GND  98.3826E-18 M=1.0 
C1500 158 162  306.8514E-18 M=1.0 
C1501 157 161  306.8514E-18 M=1.0 
C1502 152 153  55.3986E-18 M=1.0 
C1503 151 158  120.9051E-18 M=1.0 
C1504 151 157  120.9051E-18 M=1.0 
C1505 151 154  224.6967E-18 M=1.0 
C1506 151 153  224.6967E-18 M=1.0 
C1507 148 151  65.31255E-18 M=1.0 
C1508 147 152  34.9776E-18 M=1.0 
C1509 147 151  65.31255E-18 M=1.0 
C1510 OUT_2 162  55.3986E-18 M=1.0 
C1511 VDD 152  1.42083675E-15 M=1.0 
C1512 GND 162  559.068525E-18 M=1.0 
C1513 GND 161  559.068525E-18 M=1.0 
C1514 GND 158  113.0463E-18 M=1.0 
C1515 GND 157  113.0463E-18 M=1.0 
C1516 GND 151  2.3541309E-15 M=1.0 
C1517 OUT_3 161  55.3986E-18 M=1.0 
C1518 148 151  223.1748E-18 M=1.0 
C1519 147 151  223.1748E-18 M=1.0 
C1520 GND 151  2.156287725E-15 M=1.0 
C1521 GND 120  38.4993000000001E-18 M=1.0 
C1522 GND 152  69.1866E-18 M=1.0 
C1523 GND 120  1.10547E-15 M=1.0 
C1524 VDD 151  95.44635E-18 M=1.0 
C1525 VDD 120  90.3762E-18 M=1.0 
C1526 GND 152  31.6845E-18 M=1.0 
C1527 GND 120  261.0576E-18 M=1.0 
C1528 _DFF_OUT_0 DFF_OUT_1  55.3986E-18 M=1.0 
C1529 _DFF_OUT_0 DFF_OUT_0  110.7972E-18 M=1.0 
M1530 82 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1531 83 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1532 VDD GND 13 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1533 VDD GND 12 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1534 VDD GND 11 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1535 VDD GND 10 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1536 81 GND VDD VDD  TSMC18DP  L=1.17000001864653E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1537 87 86 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1538 66 65 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1539 9 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1540 93 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1541 VDD 66 93 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1542 93 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1543 84 66 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1544 VDD 86 84 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1545 84 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1546 76 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1547 VDD 65 76 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1548 76 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1549 70 86 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1550 VDD 65 70 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1551 70 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1552 28 9 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1553 VDD 86 28 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1554 28 65 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1555 16 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1556 VDD 9 16 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1557 16 65 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1558 2 66 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1559 VDD 9 2 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1560 2 86 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1561 1 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1562 VDD 66 1 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1563 1 9 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1564 91 CLK A0 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1565 71 CLK A1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1566 14 CLK A2 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1567 86 92 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1568 85 91 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1569 65 72 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1570 64 71 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1571 8 15 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1572 7 14 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1573 92 108 85 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1574 72 108 64 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1575 15 108 7 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1576 92 86 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1577 91 85 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1578 72 65 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1579 71 64 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1580 15 8 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1581 14 7 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1582 110 109 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1583 109 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1584 112 111 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1585 111 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1586 108 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1587 _DFF_OUT_0 113 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1588 _DFF_OUT_6 119 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1589 _DFF_OUT_5 118 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1590 _DFF_OUT_4 117 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1591 _DFF_OUT_3 116 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1592 _DFF_OUT_2 115 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1593 _DFF_OUT_1 114 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1594 DFF_OUT_6 _DFF_OUT_6 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1595 DFF_OUT_5 _DFF_OUT_5 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1596 DFF_OUT_4 _DFF_OUT_4 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1597 DFF_OUT_3 _DFF_OUT_3 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1598 DFF_OUT_2 _DFF_OUT_2 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1599 DFF_OUT_1 _DFF_OUT_1 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1600 DFF_OUT_0 _DFF_OUT_0 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1601 102 95 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1602 101 94 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1603 107 100 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1604 106 99 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1605 105 98 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1606 104 97 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1607 103 96 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1608 146 142 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1609 145 141 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1610 144 140 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1611 143 139 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1612 142 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1613 141 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1614 140 128 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1615 VDD 127 142 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1616 VDD 128 141 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1617 VDD 127 140 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1618 142 138 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1619 141 137 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1620 139 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1621 140 136 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1622 VDD 128 139 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1623 138 128 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1624 137 127 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1625 139 127 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1626 136 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1627 _DFF_OUT_2 _DFF_OUT_1 134 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1628 _DFF_OUT_2 _DFF_OUT_0 133 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1629 _DFF_OUT_4 _DFF_OUT_3 135 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1630 135 DFF_OUT_3 DFF_OUT_4 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1631 134 DFF_OUT_1 DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1632 133 DFF_OUT_0 DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1633 VDD 135 132 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1634 VDD 134 131 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1635 VDD 133 130 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1636 126 135 129 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1637 125 134 128 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1638 124 133 127 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1639 _DFF_OUT_6 _DFF_OUT_5 126 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1640 _DFF_OUT_6 _DFF_OUT_5 125 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1641 _DFF_OUT_6 _DFF_OUT_4 124 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1642 129 132 123 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1643 128 131 122 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1644 127 130 121 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1645 126 DFF_OUT_5 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1646 125 DFF_OUT_5 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1647 124 DFF_OUT_4 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1648 121 124 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1649 123 126 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1650 122 125 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1651 120 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1652 150 152 H_0 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1653 149 152 H_1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1654 148 152 H_2 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1655 147 152 H_3 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1656 H_1 142 DFF_OUT_4 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1657 H_1 146 _DFF_OUT_4 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1658 H_2 141 DFF_OUT_5 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1659 H_2 145 _DFF_OUT_5 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1660 H_0 140 DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1661 H_0 144 _DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1662 H_3 139 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1663 H_3 143 _DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1664 94 111 3 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1665 100 111 6 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1666 99 111 90 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1667 98 111 5 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1668 97 111 89 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1669 96 111 4 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1670 95 111 88 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1671 VDD 110 83 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1672 VDD 110 82 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1673 VDD 110 81 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1674 13 110 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1675 12 110 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1676 11 110 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1677 10 110 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1678 160 151 156 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1679 159 151 155 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1680 158 151 154 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1681 157 151 153 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1682 119 112 107 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1683 118 112 106 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1684 117 112 105 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1685 116 112 104 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1686 115 112 103 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1687 114 112 102 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1688 113 112 101 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1689 160 164 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1690 159 163 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1691 158 162 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1692 157 161 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1693 117 _DFF_OUT_4 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1694 116 _DFF_OUT_3 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1695 115 _DFF_OUT_2 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1696 114 _DFF_OUT_1 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1697 113 _DFF_OUT_0 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1698 119 _DFF_OUT_6 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1699 118 _DFF_OUT_5 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1700 99 106 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1701 98 105 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1702 97 104 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1703 96 103 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1704 95 102 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1705 94 101 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1706 100 107 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1707 OUT_0 164 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1708 OUT_1 163 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1709 OUT_2 162 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1710 OUT_3 161 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1711 162 158 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1712 161 157 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1713 164 160 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1714 163 159 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1715 156 150 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1716 155 149 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1717 154 148 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1718 153 147 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1719 152 151 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1720 151 120 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1721 90 83 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1722 89 82 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1723 88 81 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1724 VDD 13 6 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1725 VDD 12 5 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1726 VDD 11 4 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1727 VDD 10 3 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1728 86 92 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1729 85 91 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1730 65 72 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1731 64 71 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1732 8 15 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1733 7 14 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1734 87 86 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1735 66 65 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1736 9 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1737 92 86 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1738 91 85 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1739 72 65 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1740 71 64 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1741 14 7 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1742 15 8 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1743 110 109 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1744 109 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1745 91 108 A0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1746 71 108 A1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1747 14 108 A2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1748 112 111 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1749 111 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1750 108 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1751 92 CLK 85 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1752 72 CLK 64 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1753 15 CLK 7 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1754 _DFF_OUT_0 113 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1755 _DFF_OUT_6 119 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1756 _DFF_OUT_5 118 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1757 _DFF_OUT_4 117 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1758 _DFF_OUT_3 116 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1759 _DFF_OUT_2 115 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1760 _DFF_OUT_1 114 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1761 DFF_OUT_6 _DFF_OUT_6 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1762 DFF_OUT_5 _DFF_OUT_5 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1763 DFF_OUT_4 _DFF_OUT_4 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1764 DFF_OUT_3 _DFF_OUT_3 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1765 DFF_OUT_2 _DFF_OUT_2 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1766 DFF_OUT_1 _DFF_OUT_1 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1767 DFF_OUT_0 _DFF_OUT_0 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1768 105 98 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1769 104 97 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1770 103 96 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1771 102 95 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1772 101 94 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1773 107 100 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1774 106 99 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1775 142 129 189 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1776 141 129 188 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1777 189 127 187 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1778 188 128 186 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1779 140 128 185 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1780 187 138 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1781 186 137 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1782 185 127 184 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1783 184 136 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1784 139 129 183 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1785 183 128 182 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1786 182 127 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1787 93 87 181 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1788 181 66 180 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1789 180 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1790 84 66 179 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1791 179 86 178 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1792 178 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1793 76 87 177 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1794 177 65 176 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1795 176 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1796 70 86 175 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1797 175 65 174 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1798 174 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1799 28 9 173 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1800 173 86 172 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1801 172 65 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1802 16 87 171 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1803 171 9 170 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1804 170 65 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1805 2 66 169 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1806 169 9 168 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1807 168 86 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1808 1 87 167 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1809 167 66 166 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1810 166 9 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1811 150 151 H_0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1812 149 151 H_1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1813 148 151 H_2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1814 147 151 H_3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1815 H_1 146 DFF_OUT_4 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1816 H_1 142 _DFF_OUT_4 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1817 H_2 145 DFF_OUT_5 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1818 H_2 141 _DFF_OUT_5 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1819 H_0 144 DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1820 H_0 140 _DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1821 H_3 143 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1822 H_3 139 _DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1823 146 142 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1824 145 141 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1825 144 140 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1826 143 139 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1827 138 128 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1828 137 127 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1829 136 129 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1830 _DFF_OUT_2 DFF_OUT_1 134 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1831 _DFF_OUT_2 DFF_OUT_0 133 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1832 _DFF_OUT_4 DFF_OUT_3 135 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1833 135 _DFF_OUT_3 DFF_OUT_4 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1834 134 _DFF_OUT_1 DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1835 133 _DFF_OUT_0 DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1836 GND 135 132 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1837 GND 134 131 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1838 GND 133 130 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1839 126 132 129 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1840 125 131 128 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1841 124 130 127 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1842 _DFF_OUT_6 DFF_OUT_5 126 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1843 _DFF_OUT_6 DFF_OUT_5 125 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1844 _DFF_OUT_6 DFF_OUT_4 124 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1845 129 135 123 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1846 128 134 122 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1847 127 133 121 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1848 126 _DFF_OUT_5 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1849 125 _DFF_OUT_5 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1850 124 _DFF_OUT_4 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1851 121 124 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1852 123 126 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1853 122 125 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1854 120 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1855 94 112 3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1856 100 112 6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1857 99 112 90 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1858 98 112 5 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1859 97 112 89 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1860 96 112 4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1861 95 112 88 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1862 83 1 83 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1863 82 1 82 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1864 81 1 81 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1865 81 2 74 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1866 83 2 80 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1867 82 2 79 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1868 80 16 78 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1869 79 16 77 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1870 74 16 74 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1871 78 28 75 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1872 77 28 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1873 74 28 74 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1874 74 93 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1875 75 93 73 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1876 68 93 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1877 73 84 73 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1878 68 84 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1879 67 84 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1880 73 76 73 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1881 68 76 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1882 67 76 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1883 68 70 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1884 67 70 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1885 73 70 69 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1886 69 110 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1887 68 110 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1888 67 110 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1889 GND 110 63 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1890 GND 110 62 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1891 GND 110 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1892 GND 110 60 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1893 63 70 61 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1894 62 70 58 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1895 57 70 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1896 60 70 60 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1897 58 76 58 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1898 57 76 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1899 60 76 26 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1900 61 76 59 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1901 59 84 25 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1902 58 84 27 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1903 57 84 24 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1904 26 84 26 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1905 26 93 23 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1906 25 93 25 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1907 27 93 19 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1908 24 93 24 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1909 25 28 22 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1910 19 28 19 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1911 24 28 18 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1912 23 28 21 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1913 22 16 20 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1914 19 16 19 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1915 18 16 18 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1916 21 16 17 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1917 20 2 13 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1918 19 2 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1919 18 2 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1920 17 2 10 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1921 13 1 13 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1922 12 1 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1923 11 1 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1924 10 1 10 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1925 160 164 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1926 159 163 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1927 158 162 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1928 157 161 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1929 117 _DFF_OUT_4 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1930 116 _DFF_OUT_3 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1931 115 _DFF_OUT_2 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1932 114 _DFF_OUT_1 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1933 113 _DFF_OUT_0 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1934 119 _DFF_OUT_6 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1935 118 _DFF_OUT_5 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1936 99 106 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1937 98 105 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1938 97 104 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1939 96 103 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1940 95 102 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1941 94 101 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1942 100 107 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1943 OUT_0 164 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1944 OUT_1 163 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1945 OUT_2 162 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1946 OUT_3 161 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1947 162 158 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1948 161 157 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1949 164 160 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1950 163 159 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1951 160 152 156 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1952 159 152 155 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1953 158 152 154 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1954 157 152 153 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1955 156 150 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1956 155 149 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1957 154 148 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1958 153 147 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1959 152 151 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1960 151 120 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1961 119 111 107 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1962 118 111 106 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1963 117 111 105 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1964 116 111 104 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1965 115 111 103 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1966 114 111 102 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1967 113 111 101 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1968 90 83 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1969 89 82 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1970 88 81 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1971 GND 13 6 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1972 GND 12 5 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1973 GND 11 4 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1974 GND 10 3 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS PART1_G1 
 
* END OF NETLIST
.TRAN  5.00000E-11 1.50000E-08 START=  0.0000    
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
+        DELMAX = 1.00000E-10

.MEAS TRAN avg_power AVG POWER FROM=1n TO=9n
.option POST=2
.END
