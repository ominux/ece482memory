* # FILE NAME: /HOME/ENGR/TRUTY1/CADENCE/SIMULATION/WHOLE_CKT/HSPICES/          
* SCHEMATIC/NETLIST/WHOLE_CKT.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON NOV 16 12:59:16 2009
   
* GLOBAL NET DEFINITIONS
.lib "/apps/Linux/cadence-Sept2009/ncsu-cdk-1.5.1/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "/apps/Linux/cadence-Sept2009/ncsu-cdk-1.5.1/models/hspice/public/publicModel/tsmc18dN" NMOS 
.GLOBAL VDD! 
* FILE NAME: ECE482MEMORY_WHOLE_CKT_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: WHOLE_CKT.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
XI32_3 H_3 OUT_3 NET023_0 CLK_D3_ CLK_D3 REG3A_G7 
XI32_2 H_2 OUT_2 NET023_1 CLK_D3_ CLK_D3 REG3A_G7 
XI32_1 H_1 OUT_1 NET023_2 CLK_D3_ CLK_D3 REG3A_G7 
XI32_0 H_0 OUT_0 NET023_3 CLK_D3_ CLK_D3 REG3A_G7 
C0 OUT_3 0  50E-15 M=1.0 
C3 OUT_0 0  50E-15 M=1.0 
C2 OUT_1 0  50E-15 M=1.0 
C1 OUT_2 0  50E-15 M=1.0 
XI31 DFF_OUT_6 DFF_OUT_5 DFF_OUT_4 DFF_OUT_3 DFF_OUT_2 DFF_OUT_1 DFF_OUT_0 
+_DFF_OUT_6 _DFF_OUT_5 _DFF_OUT_4 _DFF_OUT_3 _DFF_OUT_2 _DFF_OUT_1 _DFF_OUT_0 
+H_0 H_1 H_2 H_3 HAMMING_7_4_G8 
XI9_6 S1OUT_6 DFF_OUT_6 _DFF_OUT_6 CLK_D2 CLK_D2_ REG2A_G9 
XI9_5 S1OUT_5 DFF_OUT_5 _DFF_OUT_5 CLK_D2 CLK_D2_ REG2A_G9 
XI9_4 S1OUT_4 DFF_OUT_4 _DFF_OUT_4 CLK_D2 CLK_D2_ REG2A_G9 
XI9_3 S1OUT_3 DFF_OUT_3 _DFF_OUT_3 CLK_D2 CLK_D2_ REG2A_G9 
XI9_2 S1OUT_2 DFF_OUT_2 _DFF_OUT_2 CLK_D2 CLK_D2_ REG2A_G9 
XI9_1 S1OUT_1 DFF_OUT_1 _DFF_OUT_1 CLK_D2 CLK_D2_ REG2A_G9 
XI9_0 S1OUT_0 DFF_OUT_0 _DFF_OUT_0 CLK_D2 CLK_D2_ REG2A_G9 
XI8 A0 A1 A2 NET051 NET050 NET049 NET048 NET047 NET046 CLK CLK_D0_ 0 VDD! 
+REG_FILE1_G10 
XI0 NET051 NET050 NET049 NET048 NET047 NET046 CLK_D1 S1OUT_6 S1OUT_5 S1OUT_4 
+S1OUT_3 S1OUT_2 S1OUT_1 S1OUT_0 0 VDD! STAGE_1_G11 
XI52 CLK NET069 INV_1 
XI59 CLK_D3_ CLK_D3 INV_2 
XI56 NET081 NET066 INV_3 
XI58 CLK_D2 CLK_D2_ INV_4 
XI49 CLK CLK_D1_ INV_5 
XI54 NET067 CLK_D3_ INV_4 
XI61 NET068 NET067 INV_5 
XI53 CLK NET068 INV_5 
XI39 CLK CLK_D0_ INV_2 
XI50 NET066 CLK_D1 INV_6 
XI51 NET069 CLK_D2 INV_7 
XI55 CLK_D1_ NET081 INV_8 
VA2_GEN A2 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 6.4E-9 12.8E-9 
V1 CLK 0  PULSE 0.0 1.8 0.0 80E-12 80E-12 700E-12 1.6E-9 
VA0_GEN A0 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 1.6E-9 3.2E-9 
VA1_GEN A1 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 3.2E-9 6.4E-9 
V0 VDD! 0  1.8 
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_8 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_8 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_4 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(810E-9) AD=+3.64500000E-13 
+AS=+3.64500000E-13 PD=+2.52000000E-06 PS=+2.52000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_4 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_3 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_3 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(450E-9) AD=+2.02500000E-13 
+AS=+2.02500000E-13 PD=+1.80000000E-06 PS=+1.80000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(900E-9) AD=+4.05000000E-13 
+AS=+4.05000000E-13 PD=+2.70000000E-06 PS=+2.70000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(630E-9) AD=+2.83500000E-13 
+AS=+2.83500000E-13 PD=+2.16000000E-06 PS=+2.16000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_6 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_6 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_7 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(630E-9) AD=+2.83500000E-13 
+AS=+2.83500000E-13 PD=+2.16000000E-06 PS=+2.16000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_7 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_5 A Y 
M0 Y A 0 0  TSMC18DN  L=(270E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(270E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_5 
   
   
   
* FILE NAME: ECE482MEMORY_NAND3_1X_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NAND3_1X.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: A<2> = A_2
*                   A<1> = A_1
*                   A<0> = A_0
*                   DOUT_ = DOUT_
*                   GND = GND
*                   VDD = VDD
.SUBCKT NAND3_1X_G3 A_2 A_1 A_0 DOUT_ GND VDD 
MP3 DOUT_ A_1 VDD VDD  TSMC18DP  L=180E-9 W=540E-9 AD=243E-15 AS=243E-15 
+PD=1.98E-6 PS=1.98E-6 M=1 
MP4 DOUT_ A_2 VDD VDD  TSMC18DP  L=180E-9 W=540E-9 AD=243E-15 AS=243E-15 
+PD=1.98E-6 PS=1.98E-6 M=1 
MP5 DOUT_ A_0 VDD VDD  TSMC18DP  L=180E-9 W=540E-9 AD=243E-15 AS=243E-15 
+PD=1.98E-6 PS=1.98E-6 M=1 
MN5 NET0111 A_1 NET0115 GND  TSMC18DN  L=180E-9 W=810E-9 AD=364.5E-15 
+AS=364.5E-15 PD=2.52E-6 PS=2.52E-6 M=1 
MN4 NET0115 A_2 GND GND  TSMC18DN  L=180E-9 W=810E-9 AD=364.5E-15 AS=364.5E-15 
+PD=2.52E-6 PS=2.52E-6 M=1 
MN6 DOUT_ A_0 NET0111 GND  TSMC18DN  L=180E-9 W=810E-9 AD=364.5E-15 
+AS=364.5E-15 PD=2.52E-6 PS=2.52E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND3_1X_G3 
* FILE NAME: ECE482MEMORY_T-GATE2_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: T-GATE2.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
*                   GND = GND
*                   PASS = PASS
*                   PASS_BAR = PASS_BAR
*                   VDD = VDD
.SUBCKT SUB1 IN OUT GND PASS PASS_BAR VDD 
M0 OUT PASS_BAR IN VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1 OUT PASS IN GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
C2 VDD PASS_BAR  26.7138E-18 M=1.0 
C3 GND PASS_BAR  21.2139E-18 M=1.0 
C4 GND PASS  43.2135E-18 M=1.0 
C5 OUT PASS_BAR  62.3646E-18 M=1.0 
C6 OUT PASS  62.3646E-18 M=1.0 
C7 GND OUT  38.5506E-18 M=1.0 
C8 IN VDD  27.1404E-18 M=1.0 
C9 IN GND  46.1574E-18 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB1 
* FILE NAME: ECE482MEMORY_REG3A_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: REG3A.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: D = D
*                   Q = Q
*                   Q_BAR = Q_BAR
*                   CLK_ = CLK_
*                   CLK = CLK
.SUBCKT REG3A_G7 D Q Q_BAR CLK_ CLK 
XI40 NODE3 0 Q_BAR VDD! INV3_G1 
XI61 NODE1 0 NODE2 VDD! INV3_G1 
XI64 NODE2 NODE3 0 CLK CLK_ VDD! SUB1 
XI63 NET27 NODE1 0 CLK_ CLK VDD! SUB2 
XI67 D 0 NET27 VDD! INV2_G2 
XI54 Q_BAR 0 Q VDD! INV2_G2 
XI55 NODE2 0 NODE1 VDD! SUB3 
XI57 Q_BAR 0 NODE3 VDD! SUB3 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS REG3A_G7 
* FILE NAME: ECE482MEMORY_REG2A_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: REG2A.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: D = D
*                   Q = Q
*                   Q_BAR = Q_BAR
*                   CLK_ = CLK_
*                   CLK = CLK
.SUBCKT REG2A_G9 D Q Q_BAR CLK_ CLK 
XI63 REG_IN NODE1 0 CLK_ CLK VDD! SUB2 
XI40 NODE3 0 Q_BAR VDD! INV3_G1 
XI61 NODE1 0 NODE2 VDD! INV3_G1 
XI64 NODE2 NODE3 0 CLK CLK_ VDD! SUB1 
XI66 D 0 REG_IN VDD! INV2_G2 
XI54 Q_BAR 0 Q VDD! INV2_G2 
XI55 NODE2 0 NODE1 VDD! SUB3 
XI57 Q_BAR 0 NODE3 VDD! SUB3 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS REG2A_G9 
* FILE NAME: ECE482MEMORY_INV0.25_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: INV0.25.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: IN = IN
*                   GND = GND
*                   OUT = OUT
*                   VDD = VDD
.SUBCKT SUB3 IN GND OUT VDD 
M0 OUT IN VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1 OUT IN GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
C2 IN VDD  26.7138E-18 M=1.0 
C3 IN GND  97.4268E-18 M=1.0 
C4 OUT VDD  27.1404E-18 M=1.0 
C5 OUT GND  84.1914E-18 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB3 
* FILE NAME: ECE482MEMORY_INV_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
.SUBCKT INV_G4 IN OUT 
MN2 OUT IN 0 0  TSMC18DN  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
MP1 OUT IN VDD! VDD!  TSMC18DP  L=180E-9 W=540E-9 AD=243E-15 AS=243E-15 
+PD=1.98E-6 PS=1.98E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_G4 
* FILE NAME: ECE482MEMORY_MUX21_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: MUX21.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   OUT = OUT
*                   SEL = SEL
*                   GND = GND
*                   VDD = VDD
.SUBCKT MUX21_G5 A B OUT SEL GND VDD 
MP2 NET13 SEL VDD VDD  TSMC18DP  L=180E-9 W=360E-9 AD=162E-15 AS=162E-15 
+PD=1.62E-6 PS=1.62E-6 M=1 
MP1 OUT SEL B VDD  TSMC18DP  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
MP0 OUT NET13 A VDD  TSMC18DP  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
MN2 NET13 SEL GND GND  TSMC18DN  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
MN1 OUT NET13 B GND  TSMC18DN  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
MN0 OUT SEL A GND  TSMC18DN  L=180E-9 W=270E-9 AD=121.5E-15 AS=121.5E-15 
+PD=1.44E-6 PS=1.44E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS MUX21_G5 
* FILE NAME: ECE482MEMORY_STAGE_1_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: STAGE_1.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A0 = A0
*                   A0_ = A0_
*                   A1 = A1
*                   A1_ = A1_
*                   A2 = A2
*                   A2_ = A2_
*                   CLK = CLK
*                   OUT<6> = OUT_6
*                   OUT<5> = OUT_5
*                   OUT<4> = OUT_4
*                   OUT<3> = OUT_3
*                   OUT<2> = OUT_2
*                   OUT<1> = OUT_1
*                   OUT<0> = OUT_0
*                   GND = GND
*                   VDD = VDD
.SUBCKT STAGE_1_G11 A0 A0_ A1 A1_ A2 A2_ CLK OUT_6 OUT_5 OUT_4 OUT_3 OUT_2 
+OUT_1 OUT_0 GND VDD 
C69 VDD A2  91.1412E-18 M=1.0 
C70 VDD A1  72.2844E-18 M=1.0 
C71 VDD A0  62.856E-18 M=1.0 
C72 A2_ VDD  62.856E-18 M=1.0 
C73 A1_ VDD  53.4276000000001E-18 M=1.0 
C74 GND 52  230.9958E-18 M=1.0 
C75 GND 51  318.9942E-18 M=1.0 
C76 GND 46  230.9958E-18 M=1.0 
C77 GND 39  324.4941E-18 M=1.0 
C78 GND 13  318.9942E-18 M=1.0 
C79 GND 3  230.9958E-18 M=1.0 
C80 GND 2  307.9944E-18 M=1.0 
C81 GND 1  230.9958E-18 M=1.0 
C82 GND A2  128.8548E-18 M=1.0 
C83 GND A1  128.8548E-18 M=1.0 
C84 GND A0  147.7116E-18 M=1.0 
C85 GND VDD  958.161149999997E-18 M=1.0 
C86 GND A2_  147.7116E-18 M=1.0 
C87 GND A1_  166.5684E-18 M=1.0 
C88 A0_ VDD  53.4276000000001E-18 M=1.0 
C89 A0_ GND  204.282E-18 M=1.0 
C90 CLK VDD  236.4957E-18 M=1.0 
C91 CLK GND  370.0647E-18 M=1.0 
C92 43 51  62.3646E-18 M=1.0 
C93 43 46  62.3646E-18 M=1.0 
C94 41 52  62.3646E-18 M=1.0 
C95 41 51  62.3646E-18 M=1.0 
C96 41 46  62.3646E-18 M=1.0 
C97 40 51  62.3646E-18 M=1.0 
C98 40 46  62.3646E-18 M=1.0 
C99 39 41  62.3646E-18 M=1.0 
C100 39 40  62.3646E-18 M=1.0 
C101 35 39  62.3646E-18 M=1.0 
C102 33 46  62.3646E-18 M=1.0 
C103 16 46  62.3646E-18 M=1.0 
C104 16 39  62.3646E-18 M=1.0 
C105 14 51  62.3646E-18 M=1.0 
C106 13 44  62.3646E-18 M=1.0 
C107 12 52  62.3646E-18 M=1.0 
C108 11 52  62.3646E-18 M=1.0 
C109 6 13  62.3646E-18 M=1.0 
C110 3 44  62.3646E-18 M=1.0 
C111 3 6  62.3646E-18 M=1.0 
C112 3 5  62.3646E-18 M=1.0 
C113 A1 46  62.3646E-18 M=1.0 
C114 A1 39  62.3646E-18 M=1.0 
C115 A0 51  62.3646E-18 M=1.0 
C116 A0 39  124.7292E-18 M=1.0 
C117 A0 13  62.3646E-18 M=1.0 
C118 OUT_2 1  62.3646E-18 M=1.0 
C119 VDD 52  76.068E-18 M=1.0 
C120 VDD 51  76.068E-18 M=1.0 
C121 VDD 46  76.068E-18 M=1.0 
C122 VDD 39  76.068E-18 M=1.0 
C123 VDD 13  76.068E-18 M=1.0 
C124 VDD 3  76.068E-18 M=1.0 
C125 VDD 2  76.068E-18 M=1.0 
C126 VDD 1  76.068E-18 M=1.0 
C127 VDD A2  32.4936E-18 M=1.0 
C128 VDD OUT_2  63.8441999999999E-18 M=1.0 
C129 A2_ 13  124.7292E-18 M=1.0 
C130 A2_ 3  62.3646E-18 M=1.0 
C131 A2_ 2  62.3646E-18 M=1.0 
C132 OUT_1 1  62.3646E-18 M=1.0 
C133 OUT_1 VDD  63.8442E-18 M=1.0 
C134 A1_ 52  62.3646E-18 M=1.0 
C135 A1_ 51  124.7292E-18 M=1.0 
C136 A1_ 2  124.7292E-18 M=1.0 
C137 A1_ 1  62.3646E-18 M=1.0 
C138 OUT_0 1  62.3646E-18 M=1.0 
C139 OUT_0 VDD  63.8442E-18 M=1.0 
C140 GND 52  478.337399999999E-18 M=1.0 
C141 GND 51  442.683E-18 M=1.0 
C142 GND 46  349.0218E-18 M=1.0 
C143 GND 39  231.26985E-18 M=1.0 
C144 GND 13  564.391799999999E-18 M=1.0 
C145 GND 3  601.947900000001E-18 M=1.0 
C146 GND 2  757.5786E-18 M=1.0 
C147 GND 1  741.343500000001E-18 M=1.0 
C148 GND A2  571.0374E-18 M=1.0 
C149 GND A1  993.0168E-18 M=1.0 
C150 GND A0  1.1522979E-15 M=1.0 
C151 GND OUT_2  128.4579E-18 M=1.0 
C152 GND VDD  2.2258791E-15 M=1.0 
C153 GND A2_  768.1545E-18 M=1.0 
C154 GND OUT_1  128.4579E-18 M=1.0 
C155 GND A1_  1.3039722E-15 M=1.0 
C156 GND OUT_0  128.4579E-18 M=1.0 
C157 A0_ 52  124.7292E-18 M=1.0 
C158 A0_ 46  124.7292E-18 M=1.0 
C159 A0_ 3  124.7292E-18 M=1.0 
C160 A0_ 1  124.7292E-18 M=1.0 
C161 A0_ GND  1.371708E-15 M=1.0 
C162 CLK VDD  509.6133E-18 M=1.0 
C163 CLK GND  1.5018732E-15 M=1.0 
C164 OUT_6 1  62.3646E-18 M=1.0 
C165 OUT_6 VDD  63.8442E-18 M=1.0 
C166 OUT_6 GND  128.4579E-18 M=1.0 
C167 OUT_5 1  62.3646E-18 M=1.0 
C168 OUT_5 VDD  63.8442000000001E-18 M=1.0 
C169 OUT_5 GND  128.4579E-18 M=1.0 
C170 OUT_4 1  62.3646E-18 M=1.0 
C171 OUT_4 VDD  63.8442000000001E-18 M=1.0 
C172 OUT_4 GND  128.4579E-18 M=1.0 
C173 OUT_3 1  62.3646E-18 M=1.0 
C174 OUT_3 VDD  63.8441999999999E-18 M=1.0 
C175 OUT_3 GND  128.4579E-18 M=1.0 
C176 51 52  110.7972E-18 M=1.0 
C177 46 52  110.7972E-18 M=1.0 
C178 46 51  110.7972E-18 M=1.0 
C179 41 52  65.0448E-18 M=1.0 
C180 41 51  65.0448E-18 M=1.0 
C181 41 46  65.0448E-18 M=1.0 
C182 40 52  65.0448E-18 M=1.0 
C183 40 51  65.0448E-18 M=1.0 
C184 40 46  65.0448E-18 M=1.0 
C185 39 52  55.3986E-18 M=1.0 
C186 39 51  55.3986E-18 M=1.0 
C187 39 46  55.3986E-18 M=1.0 
C188 39 41  65.0448E-18 M=1.0 
C189 39 40  65.0448E-18 M=1.0 
C190 38 39  65.0448E-18 M=1.0 
C191 37 39  65.0448E-18 M=1.0 
C192 36 46  65.0448E-18 M=1.0 
C193 35 46  65.0448E-18 M=1.0 
C194 35 39  65.0448E-18 M=1.0 
C195 34 51  65.0448E-18 M=1.0 
C196 33 51  65.0448E-18 M=1.0 
C197 33 46  65.0448E-18 M=1.0 
C198 16 51  65.0448E-18 M=1.0 
C199 16 46  65.0448E-18 M=1.0 
C200 16 39  65.0448E-18 M=1.0 
C201 15 52  65.0448E-18 M=1.0 
C202 14 52  65.0448E-18 M=1.0 
C203 14 51  65.0448E-18 M=1.0 
C204 13 52  110.7972E-18 M=1.0 
C205 13 51  110.7972E-18 M=1.0 
C206 13 46  110.7972E-18 M=1.0 
C207 13 44  65.0448E-18 M=1.0 
C208 13 41  65.0448E-18 M=1.0 
C209 13 39  55.3986E-18 M=1.0 
C210 12 52  65.0448E-18 M=1.0 
C211 12 13  65.0448E-18 M=1.0 
C212 11 52  65.0448E-18 M=1.0 
C213 11 13  65.0448E-18 M=1.0 
C214 10 13  65.0448E-18 M=1.0 
C215 6 13  65.0448E-18 M=1.0 
C216 3 52  110.7972E-18 M=1.0 
C217 3 51  110.7972E-18 M=1.0 
C218 3 47  60.31485E-18 M=1.0 
C219 3 46  110.7972E-18 M=1.0 
C220 3 44  64.945575E-18 M=1.0 
C221 3 39  55.3986E-18 M=1.0 
C222 3 13  110.7972E-18 M=1.0 
C223 3 9  65.0448E-18 M=1.0 
C224 3 8  65.0448E-18 M=1.0 
C225 3 6  65.0448E-18 M=1.0 
C226 3 5  65.0448E-18 M=1.0 
C227 2 52  110.7972E-18 M=1.0 
C228 2 51  110.7972E-18 M=1.0 
C229 2 49  60.31485E-18 M=1.0 
C230 2 46  110.7972E-18 M=1.0 
C231 2 44  60.31485E-18 M=1.0 
C232 2 39  55.3986E-18 M=1.0 
C233 2 13  110.7972E-18 M=1.0 
C234 2 7  60.31485E-18 M=1.0 
C235 2 6  60.31485E-18 M=1.0 
C236 2 5  60.31485E-18 M=1.0 
C237 2 4  60.31485E-18 M=1.0 
C238 2 3  110.7972E-18 M=1.0 
C239 1 52  110.7972E-18 M=1.0 
C240 1 51  110.7972E-18 M=1.0 
C241 1 46  110.7972E-18 M=1.0 
C242 1 39  55.3986E-18 M=1.0 
C243 1 13  110.7972E-18 M=1.0 
C244 1 3  110.7972E-18 M=1.0 
C245 1 2  110.7972E-18 M=1.0 
C246 A2 51  55.3986E-18 M=1.0 
C247 A2 46  55.3986E-18 M=1.0 
C248 A2 39  55.3986E-18 M=1.0 
C249 A1 46  55.93725E-18 M=1.0 
C250 A1 39  55.93725E-18 M=1.0 
C251 A0 51  55.93725E-18 M=1.0 
C252 A0 13  55.93725E-18 M=1.0 
C253 A0 A1  221.5944E-18 M=1.0 
C254 OUT_2 1  120.70665E-18 M=1.0 
C255 VDD 52  1.3095432E-15 M=1.0 
C256 VDD 51  260.1792E-18 M=1.0 
C257 VDD 46  260.1792E-18 M=1.0 
C258 VDD 39  195.1344E-18 M=1.0 
C259 VDD 13  1.6542396E-15 M=1.0 
C260 VDD 3  874.9422E-18 M=1.0 
C261 VDD 2  874.9422E-18 M=1.0 
C262 VDD 1  1.02615435E-15 M=1.0 
C263 VDD A1  1.0080801E-15 M=1.0 
C264 VDD A0  1.0389987E-15 M=1.0 
C265 A2_ 13  55.3986E-18 M=1.0 
C266 A2_ 3  55.3986E-18 M=1.0 
C267 A2_ 2  55.3986E-18 M=1.0 
C268 A2_ 1  55.3986E-18 M=1.0 
C269 A2_ VDD  69.8679E-18 M=1.0 
C270 OUT_1 1  120.3381E-18 M=1.0 
C271 A1_ 51  55.3986E-18 M=1.0 
C272 A1_ 46  55.3986E-18 M=1.0 
C273 A1_ 39  55.3986E-18 M=1.0 
C274 A1_ 13  55.3986E-18 M=1.0 
C275 A1_ 3  55.3986E-18 M=1.0 
C276 A1_ 2  55.3986E-18 M=1.0 
C277 A1_ 1  55.3986E-18 M=1.0 
C278 A1_ A2  221.5944E-18 M=1.0 
C279 A1_ VDD  69.8679E-18 M=1.0 
C280 A1_ A2_  221.5944E-18 M=1.0 
C281 OUT_0 1  120.70665E-18 M=1.0 
C282 GND 52  5.1312726E-15 M=1.0 
C283 GND 51  4.36871205E-15 M=1.0 
C284 GND 46  4.32981045E-15 M=1.0 
C285 GND 39  3.57453E-15 M=1.0 
C286 GND 13  2.6428122E-15 M=1.0 
C287 GND 3  3.52900575E-15 M=1.0 
C288 GND 2  3.60116685E-15 M=1.0 
C289 GND 1  3.359115E-15 M=1.0 
C290 GND A2  2.1029508E-15 M=1.0 
C291 GND A1  702.2196E-18 M=1.0 
C292 GND A0  315.4158E-18 M=1.0 
C293 GND VDD  2.50304535E-15 M=1.0 
C294 GND A2_  1.4247936E-15 M=1.0 
C295 GND A1_  1.1145366E-15 M=1.0 
C296 A0_ A1  221.5944E-18 M=1.0 
C297 A0_ A0  166.1958E-18 M=1.0 
C298 A0_ VDD  1.3209156E-15 M=1.0 
C299 A0_ GND  636.5178E-18 M=1.0 
C300 CLK 1  582.5736E-18 M=1.0 
C301 CLK VDD  1.4428683E-15 M=1.0 
C302 CLK GND  7.01162145E-15 M=1.0 
C303 OUT_6 1  64.84635E-18 M=1.0 
C304 OUT_5 1  55.62945E-18 M=1.0 
C305 OUT_4 1  120.70665E-18 M=1.0 
C306 OUT_3 1  120.3381E-18 M=1.0 
M307 OUT_5 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M308 OUT_3 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M309 VDD GND OUT_6 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M310 VDD GND OUT_4 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M311 VDD GND OUT_2 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M312 VDD GND OUT_0 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M313 OUT_1 GND VDD VDD  TSMC18DP  L=1.17000001864653E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M314 VDD CLK OUT_1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M315 VDD CLK OUT_5 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M316 VDD CLK OUT_3 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M317 OUT_6 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M318 OUT_4 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M319 OUT_2 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M320 OUT_0 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M321 52 A0_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M322 VDD A1_ 52 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M323 52 A2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M324 51 A1_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M325 VDD A0 51 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M326 51 A2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M327 46 A0_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M328 VDD A1 46 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M329 46 A2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M330 39 A0 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M331 VDD A1 39 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M332 39 A2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M333 13 A2_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M334 VDD A0 13 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M335 13 A1 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M336 3 A0_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M337 VDD A2_ 3 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M338 3 A1 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M339 2 A1_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M340 VDD A2_ 2 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M341 2 A0 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M342 1 A0_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M343 VDD A1_ 1 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M344 1 A2_ VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M345 OUT_5 1 OUT_5 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M346 OUT_3 1 OUT_3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M347 OUT_1 1 OUT_1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M348 OUT_5 2 50 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M349 OUT_3 2 49 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M350 OUT_1 2 44 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M351 44 3 44 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M352 50 3 48 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M353 49 3 47 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M354 48 13 45 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M355 47 13 41 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M356 44 13 44 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M357 45 52 43 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M358 41 52 41 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M359 44 52 40 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M360 41 51 41 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M361 40 51 40 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M362 43 51 43 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M363 43 46 43 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M364 41 46 41 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M365 40 46 40 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M366 43 39 42 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M367 41 39 41 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M368 40 39 40 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M369 42 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M370 41 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M371 40 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M372 GND CLK 38 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M373 GND CLK 37 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M374 GND CLK 16 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M375 GND CLK 35 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M376 38 39 36 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M377 37 39 33 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M378 16 39 16 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M379 35 39 35 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M380 36 46 34 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M381 33 46 33 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M382 16 46 16 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M383 35 46 14 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M384 34 51 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M385 33 51 15 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M386 16 51 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M387 14 51 14 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M388 14 52 10 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M389 12 52 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M390 15 52 6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M391 11 52 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M392 12 13 9 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M393 6 13 6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M394 11 13 5 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M395 10 13 8 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M396 8 3 4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M397 9 3 7 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M398 6 3 6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M399 5 3 5 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M400 7 2 OUT_6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M401 6 2 OUT_4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M402 5 2 OUT_2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M403 4 2 OUT_0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M404 OUT_6 1 OUT_6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M405 OUT_4 1 OUT_4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M406 OUT_2 1 OUT_2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M407 OUT_0 1 OUT_0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M408 52 A0_ 68 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M409 68 A1_ 67 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M410 67 A2 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M411 51 A1_ 66 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M412 66 A0 65 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M413 65 A2 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M414 46 A0_ 64 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M415 64 A1 63 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M416 63 A2 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M417 39 A0 62 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M418 62 A1 61 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M419 61 A2 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M420 13 A2_ 60 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M421 60 A0 59 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M422 59 A1 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M423 3 A0_ 58 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M424 58 A2_ 57 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M425 57 A1 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M426 2 A1_ 56 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M427 56 A2_ 55 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M428 55 A0 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M429 1 A0_ 54 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M430 54 A1_ 53 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M431 53 A2_ GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS STAGE_1_G11 
* FILE NAME: ECE482MEMORY_HAMMING_7_4_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: HAMMING_7_4.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: B<6> = B_6
*                   B<5> = B_5
*                   B<4> = B_4
*                   B<3> = B_3
*                   B<2> = B_2
*                   B<1> = B_1
*                   B<0> = B_0
*                   B_<6> = B__6
*                   B_<5> = B__5
*                   B_<4> = B__4
*                   B_<3> = B__3
*                   B_<2> = B__2
*                   B_<1> = B__1
*                   B_<0> = B__0
*                   C0 = C0
*                   C1 = C1
*                   C2 = C2
*                   C3 = C3
.SUBCKT HAMMING_7_4_G8 B_6 B_5 B_4 B_3 B_2 B_1 B_0 B__6 B__5 B__4 B__3 B__2 
+B__1 B__0 C0 C1 C2 C3 
XI14 P0 P1 P2 NET22 0 VDD! NAND3_1X_G3 
XI15 P0_ P1 P2 NET26 0 VDD! NAND3_1X_G3 
XI16 P0 P1_ P2 NET30 0 VDD! NAND3_1X_G3 
XI17 P0 P1 P2_ NET34 0 VDD! NAND3_1X_G3 
XI13 P2 P2_ INV_G4 
XI12 P1 P1_ INV_G4 
XI11 P0 P0_ INV_G4 
XI6 B_2 B__2 C0 NET34 0 VDD! MUX21_G5 
XI5 B_4 B__4 C1 NET30 0 VDD! MUX21_G5 
XI4 B_5 B__5 C2 NET26 0 VDD! MUX21_G5 
XI3 B_6 B__6 C3 NET22 0 VDD! MUX21_G5 
XI1 B_6 B__6 B_5 B__5 B_2 B__2 B_1 B__1 P1 0 VDD! XOR4_G6 
XI0 B_6 B__6 B_4 B__4 B_2 B__2 B_0 B__0 P0 0 VDD! XOR4_G6 
XI2 B_6 B__6 B_5 B__5 B_4 B__4 B_3 B__3 P2 0 VDD! XOR4_G6 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS HAMMING_7_4_G8 
* FILE NAME: ECE482MEMORY_INV3_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: INV3.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: IN = IN
*                   GND = GND
*                   OUT = OUT
*                   VDD = VDD
.SUBCKT INV3_G1 IN GND OUT VDD 
M0 OUT IN VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1 OUT IN GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
C2 IN GND  39.285E-18 M=1.0 
C3 GND VDD  40.9689E-18 M=1.0 
C4 OUT VDD  27.1404E-18 M=1.0 
C5 OUT GND  59.4693E-18 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV3_G1 
* FILE NAME: ECE482MEMORY_INV2_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: INV2.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: IN = IN
*                   GND = GND
*                   OUT = OUT
*                   VDD = VDD
.SUBCKT INV2_G2 IN GND OUT VDD 
M0 OUT IN VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1 OUT IN GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
C2 IN GND  38.4993E-18 M=1.0 
C3 GND VDD  37.1655E-18 M=1.0 
C4 OUT VDD  27.1404E-18 M=1.0 
C5 OUT GND  67.5927E-18 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV2_G2 
* FILE NAME: ECE482MEMORY_REG_FILE1_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: REG_FILE1.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   Q0 = Q0
*                   Q0_BAR = Q0_BAR
*                   Q1 = Q1
*                   Q1_BAR = Q1_BAR
*                   Q2 = Q2
*                   Q2_BAR = Q2_BAR
*                   CLK = CLK
*                   CLK_BAR = CLK_BAR
*                   GND = GND
*                   VDD = VDD
.SUBCKT REG_FILE1_G10 D0 D1 D2 Q0 Q0_BAR Q1 Q1_BAR Q2 Q2_BAR CLK CLK_BAR GND 
+VDD 
C10 VDD 6  53.4276E-18 M=1.0 
C11 VDD 5  53.4276E-18 M=1.0 
C12 VDD 4  53.4276E-18 M=1.0 
C13 Q2 VDD  66.7845E-18 M=1.0 
C14 Q1 VDD  66.7845E-18 M=1.0 
C15 Q0 VDD  66.7845E-18 M=1.0 
C16 CLK_BAR VDD  108.4266E-18 M=1.0 
C17 GND 9  29.8566E-18 M=1.0 
C18 GND 8  29.8566E-18 M=1.0 
C19 GND 7  29.8566E-18 M=1.0 
C20 GND 6  182.2824E-18 M=1.0 
C21 GND 5  182.2824E-18 M=1.0 
C22 GND 4  182.2824E-18 M=1.0 
C23 GND 3  29.8566E-18 M=1.0 
C24 GND 2  29.8566E-18 M=1.0 
C25 GND 1  29.8566E-18 M=1.0 
C26 GND Q2  221.5674E-18 M=1.0 
C27 GND Q1  221.5674E-18 M=1.0 
C28 GND Q0  221.5674E-18 M=1.0 
C29 GND CLK_BAR  129.6405E-18 M=1.0 
C30 CLK VDD  160.2828E-18 M=1.0 
C31 CLK GND  96.6411E-18 M=1.0 
C32 VDD 9  46.674E-18 M=1.0 
C33 VDD 8  46.674E-18 M=1.0 
C34 VDD 7  46.674E-18 M=1.0 
C35 VDD 6  54.2808E-18 M=1.0 
C36 VDD 5  54.2808E-18 M=1.0 
C37 VDD 4  54.2808E-18 M=1.0 
C38 VDD 3  46.674E-18 M=1.0 
C39 VDD 2  46.674E-18 M=1.0 
C40 VDD 1  46.674E-18 M=1.0 
C41 VDD Q0_BAR  27.1404E-18 M=1.0 
C42 Q2 VDD  27.1404E-18 M=1.0 
C43 Q1 VDD  27.1404E-18 M=1.0 
C44 Q0 VDD  27.1404E-18 M=1.0 
C45 Q1_BAR VDD  27.1404E-18 M=1.0 
C46 CLK_BAR 9  62.3646E-18 M=1.0 
C47 CLK_BAR 8  62.3646E-18 M=1.0 
C48 CLK_BAR 7  62.3646E-18 M=1.0 
C49 CLK_BAR 3  62.3646E-18 M=1.0 
C50 CLK_BAR 2  62.3646E-18 M=1.0 
C51 CLK_BAR 1  62.3646E-18 M=1.0 
C52 CLK_BAR VDD  53.5221E-18 M=1.0 
C53 GND 9  205.6968E-18 M=1.0 
C54 GND 8  205.6968E-18 M=1.0 
C55 GND 7  205.6968E-18 M=1.0 
C56 GND 6  167.6628E-18 M=1.0 
C57 GND 5  167.6628E-18 M=1.0 
C58 GND 4  167.6628E-18 M=1.0 
C59 GND 3  188.6859E-18 M=1.0 
C60 GND 2  188.6859E-18 M=1.0 
C61 GND 1  188.6859E-18 M=1.0 
C62 GND Q0_BAR  93.6999E-18 M=1.0 
C63 GND VDD  984.6612E-18 M=1.0 
C64 GND Q2  172.2303E-18 M=1.0 
C65 GND Q1  172.2303E-18 M=1.0 
C66 GND Q0  172.2303E-18 M=1.0 
C67 GND Q1_BAR  93.6999E-18 M=1.0 
C68 GND CLK_BAR  127.2591E-18 M=1.0 
C69 Q2_BAR VDD  27.1404E-18 M=1.0 
C70 Q2_BAR GND  93.6999E-18 M=1.0 
C71 CLK 6  62.3646E-18 M=1.0 
C72 CLK 5  62.3646E-18 M=1.0 
C73 CLK 4  62.3646E-18 M=1.0 
C74 CLK 3  62.3646E-18 M=1.0 
C75 CLK 2  62.3646E-18 M=1.0 
C76 CLK 1  62.3646E-18 M=1.0 
C77 CLK VDD  127.0944E-18 M=1.0 
C78 D2 VDD  27.1404E-18 M=1.0 
C79 D2 GND  74.6829E-18 M=1.0 
C80 D1 VDD  27.1404E-18 M=1.0 
C81 D1 GND  65.1744E-18 M=1.0 
C82 D0 VDD  27.1404E-18 M=1.0 
C83 D0 GND  76.5846E-18 M=1.0 
C84 3 6  342.873E-18 M=1.0 
C85 2 5  342.873E-18 M=1.0 
C86 1 4  342.873E-18 M=1.0 
C87 VDD 9  34.9776E-18 M=1.0 
C88 VDD 8  34.9776E-18 M=1.0 
C89 VDD 7  34.9776E-18 M=1.0 
C90 VDD 6  65.5065E-18 M=1.0 
C91 VDD 5  65.5065E-18 M=1.0 
C92 VDD 4  65.5065E-18 M=1.0 
C93 VDD 3  34.9776E-18 M=1.0 
C94 VDD 2  34.9776E-18 M=1.0 
C95 VDD 1  34.9776E-18 M=1.0 
C96 Q2 9  345.2904E-18 M=1.0 
C97 Q2 VDD  65.5065E-18 M=1.0 
C98 Q1 8  345.2904E-18 M=1.0 
C99 Q1 VDD  65.5065E-18 M=1.0 
C100 Q0 7  345.2904E-18 M=1.0 
C101 Q0 Q0_BAR  55.3986E-18 M=1.0 
C102 Q0 VDD  65.5065E-18 M=1.0 
C103 Q1_BAR Q1  55.3986E-18 M=1.0 
C104 CLK_BAR 9  55.3986E-18 M=1.0 
C105 CLK_BAR 8  55.3986E-18 M=1.0 
C106 CLK_BAR 7  55.3986E-18 M=1.0 
C107 CLK_BAR 6  201.6873E-18 M=1.0 
C108 CLK_BAR 5  201.6873E-18 M=1.0 
C109 CLK_BAR 4  201.6873E-18 M=1.0 
C110 CLK_BAR 3  75.29535E-18 M=1.0 
C111 CLK_BAR 2  75.29535E-18 M=1.0 
C112 CLK_BAR 1  75.29535E-18 M=1.0 
C113 GND 9  57.4344E-18 M=1.0 
C114 GND 8  57.4344E-18 M=1.0 
C115 GND 7  57.4344E-18 M=1.0 
C116 GND 6  222.9867E-18 M=1.0 
C117 GND 5  222.9867E-18 M=1.0 
C118 GND 4  222.9867E-18 M=1.0 
C119 GND 3  49.167E-18 M=1.0 
C120 GND 2  49.167E-18 M=1.0 
C121 GND 1  49.167E-18 M=1.0 
C122 GND VDD  4.1364711E-15 M=1.0 
C123 GND Q2  391.5135E-18 M=1.0 
C124 GND Q1  391.5135E-18 M=1.0 
C125 GND Q0  391.5135E-18 M=1.0 
C126 GND CLK_BAR  2.77924995E-15 M=1.0 
C127 Q2_BAR Q2  55.3986E-18 M=1.0 
C128 CLK 6  143.21295E-18 M=1.0 
C129 CLK 5  143.21295E-18 M=1.0 
C130 CLK 4  143.21295E-18 M=1.0 
C131 CLK 3  90.3762E-18 M=1.0 
C132 CLK 2  90.3762E-18 M=1.0 
C133 CLK 1  90.3762E-18 M=1.0 
C134 CLK VDD  1.29330675E-15 M=1.0 
C135 D1 VDD  55.3986E-18 M=1.0 
C136 D0 VDD  55.3986E-18 M=1.0 
C137 CLK_BAR 6  69.4476E-18 M=1.0 
C138 CLK_BAR 5  69.4476E-18 M=1.0 
C139 CLK_BAR VDD  788.29965E-18 M=1.0 
C140 GND CLK_BAR  858.0897E-18 M=1.0 
C141 CLK 5  94.4298E-18 M=1.0 
C142 CLK 4  94.4298E-18 M=1.0 
C143 CLK 2  52.3044E-18 M=1.0 
C144 CLK 1  52.3044E-18 M=1.0 
C145 CLK VDD  599.2362E-18 M=1.0 
C146 CLK CLK_BAR  155.8836E-18 M=1.0 
C147 CLK GND  965.9169E-18 M=1.0 
M148 3 CLK D2 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M149 2 CLK D1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M150 1 CLK D0 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M151 9 CLK_BAR 6 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M152 8 CLK_BAR 5 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M153 7 CLK_BAR 4 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M154 Q2 9 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M155 Q1 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M156 Q0 7 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M157 4 1 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M158 6 3 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M159 5 2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M160 9 Q2 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M161 8 Q1 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M162 7 Q0 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M163 3 6 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M164 2 5 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M165 1 4 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M166 Q2_BAR Q2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M167 Q1_BAR Q1 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M168 Q0_BAR Q0 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M169 3 CLK_BAR D2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M170 2 CLK_BAR D1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M171 1 CLK_BAR D0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M172 9 CLK 6 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M173 8 CLK 5 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M174 7 CLK 4 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M175 Q1 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M176 Q0 7 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M177 Q2 9 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M178 6 3 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M179 5 2 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M180 4 1 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M181 9 Q2 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M182 8 Q1 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M183 7 Q0 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M184 3 6 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M185 2 5 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M186 1 4 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M187 Q2_BAR Q2 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M188 Q1_BAR Q1 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M189 Q0_BAR Q0 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS REG_FILE1_G10 
* FILE NAME: ECE482MEMORY_XOR4_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: XOR4.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:08 2009.
   
* TERMINAL MAPPING: A = A
*                   A_ = A_
*                   B = B
*                   B_ = B_
*                   C = C
*                   C_ = C_
*                   D = D
*                   D_ = D_
*                   OUT = OUT
*                   GND = GND
*                   VDD = VDD
.SUBCKT XOR4_G6 A A_ B B_ C C_ D D_ OUT GND VDD 
C5 VDD 4  47.142E-18 M=1.0 
C6 VDD 2  21.2139E-18 M=1.0 
C7 D VDD  57.945375E-18 M=1.0 
C8 GND 4  66.7845E-18 M=1.0 
C9 GND 3  57.3561E-18 M=1.0 
C10 GND 2  25.9281E-18 M=1.0 
C11 GND D_  57.3561E-18 M=1.0 
C12 GND D  59.909625E-18 M=1.0 
C13 B VDD  78.57E-18 M=1.0 
C14 B GND  36.1422E-18 M=1.0 
C15 B_ GND  52.6419E-18 M=1.0 
C16 3 4  62.3646E-18 M=1.0 
C17 2 4  62.3646E-18 M=1.0 
C18 2 3  87.1128E-18 M=1.0 
C19 VDD 4  69.4944E-18 M=1.0 
C20 VDD 2  151.3224E-18 M=1.0 
C21 VDD 1  27.1404E-18 M=1.0 
C22 D_ 4  62.3646E-18 M=1.0 
C23 OUT 3  62.3646E-18 M=1.0 
C24 OUT VDD  27.1404E-18 M=1.0 
C25 D 4  62.3646E-18 M=1.0 
C26 C VDD  36.5499E-18 M=1.0 
C27 C D_  62.3646E-18 M=1.0 
C28 GND 4  448.4826E-18 M=1.0 
C29 GND 3  39.1662E-18 M=1.0 
C30 GND 2  94.068E-18 M=1.0 
C31 GND 1  46.1574E-18 M=1.0 
C32 GND D_  20.0502E-18 M=1.0 
C33 GND OUT  51.1479E-18 M=1.0 
C34 GND D  20.0502E-18 M=1.0 
C35 GND C  38.5506E-18 M=1.0 
C36 B 2  105.67395E-18 M=1.0 
C37 A VDD  27.1404E-18 M=1.0 
C38 A GND  59.1174E-18 M=1.0 
C39 C_ VDD  27.1404E-18 M=1.0 
C40 C_ D  62.3646E-18 M=1.0 
C41 C_ GND  58.1391E-18 M=1.0 
C42 B_ 2  62.3646E-18 M=1.0 
C43 B_ GND  20.1546E-18 M=1.0 
C44 B_ A  62.3646E-18 M=1.0 
C45 A_ VDD  36.5499E-18 M=1.0 
C46 A_ GND  24.1614E-18 M=1.0 
C47 A_ B  152.442E-18 M=1.0 
C48 2 3  34.9776E-18 M=1.0 
C49 1 2  55.3986E-18 M=1.0 
C50 VDD 2  130.5198E-18 M=1.0 
C51 OUT 2  55.3986E-18 M=1.0 
C52 GND 2  74.1006E-18 M=1.0 
M53 C_ D_ 4 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M54 4 D C VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M55 VDD 4 3 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M56 2 4 OUT VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M57 A_ B_ 2 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M58 OUT 3 1 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M59 2 B A VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M60 1 2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M61 2 3 OUT GND  TSMC18DN  L=180.000000682412E-9 W=360.000001364824E-9 
+AD=161.999997834797E-15 AS=97.1999987008781E-15 PD=1.25999997635518E-6 
+PS=539.999973625527E-9 M=1 
M62 OUT 4 1 GND  TSMC18DN  L=180.000000682412E-9 W=360.000001364824E-9 
+AD=97.1999987008781E-15 AS=97.1999987008781E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M63 1 2 GND GND  TSMC18DN  L=180.000000682412E-9 W=360.000001364824E-9 
+AD=97.1999987008781E-15 AS=161.999997834797E-15 PD=539.999973625527E-9 
+PS=1.25999997635518E-6 M=1 
M64 C_ D 4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M65 4 D_ C GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M66 GND 4 3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M67 A_ B 2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M68 2 B_ A GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS XOR4_G6 
* FILE NAME: ECE482MEMORY_T-GATE_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: T-GATE.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  6 16:40:07 2009.
   
* TERMINAL MAPPING: IN = IN
*                   OUT = OUT
*                   GND = GND
*                   PASS = PASS
*                   PASS_BAR = PASS_BAR
*                   VDD = VDD
.SUBCKT SUB2 IN OUT GND PASS PASS_BAR VDD 
M0 OUT PASS_BAR IN VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1 OUT PASS IN GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
C2 VDD PASS_BAR  26.7138E-18 M=1.0 
C3 GND PASS_BAR  21.9996E-18 M=1.0 
C4 GND PASS  43.2135E-18 M=1.0 
C5 OUT PASS_BAR  62.3646E-18 M=1.0 
C6 OUT PASS  62.3646E-18 M=1.0 
C7 GND OUT  30.9438E-18 M=1.0 
C8 IN VDD  27.1404E-18 M=1.0 
C9 IN GND  38.5506E-18 M=1.0 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB2 
 
* END OF NETLIST
.TRAN  5.00000E-11 1.50000E-08 START=  0.0000    
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
+        DELMAX = 1.00000E-10

.MEAS TRAN avg_power AVG POWER FROM=1n TO=9n
.option POST=2
.END
