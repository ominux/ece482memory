* # FILE NAME: /HOME/ENGR/TRUTY1/CADENCE/SIMULATION/WHOLE_CKT/HSPICES/          
* SCHEMATIC/NETLIST/WHOLE_CKT.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON NOV 16 12:59:16 2009
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: PROJECT_WHOLE_CKT_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: WHOLE_CKT.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
.lib "/apps/Linux/cadence-Sept2009/ncsu-cdk-1.5.1/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "/apps/Linux/cadence-Sept2009/ncsu-cdk-1.5.1/models/hspice/public/publicModel/tsmc18dN" NMOS 
  
XI6 CLK NET06 INV_1 
XI7 NET06 CLK_D INV_2 
XI2 A1 A1_ INV_3 
XI1 A0 A0_ INV_3 
XI4_2 OUT_2 NET048_0 INV_1 
XI4_1 OUT_1 NET048_1 INV_1 
XI4_0 OUT_0 NET048_2 INV_1 
XI5_2 NET048_0 DFF_OUT_2 INV_4 
XI5_1 NET048_1 DFF_OUT_1 INV_4 
XI5_0 NET048_2 DFF_OUT_0 INV_4 
XI3 A2 A2_ INV_3 
XI0 A0 A0_ A1 A1_ A2 A2_ CLK_D OUT_6 OUT_5 OUT_4 OUT_3 OUT_2 OUT_1 OUT_0 0 
+VDD! STAGE_1_G4 
VA2_GEN A2 0  PULSE 1.8 0.0 80E-12 80E-12 80E-12 6.4E-9 12.8E-9 
V1 CLK 0  PULSE 0.0 1.8 0.0 80E-12 80E-12 700E-12 1.6E-9 
VA0_GEN A0 0  PULSE 1.8 0.0 80E-12 80E-12 80E-12 1.6E-9 3.2E-9 
VA1_GEN A1 0  PULSE 1.8 0.0 80E-12 80E-12 80E-12 3.2E-9 6.4E-9 
V0 VDD! 0  1.8 
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(270E-9) AD=+1.21500000E-13 
+AS=+1.21500000E-13 PD=+1.44000000E-06 PS=+1.44000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_3 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(540E-9) AD=+2.43000000E-13 
+AS=+2.43000000E-13 PD=+1.98000000E-06 PS=+1.98000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_3 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_4 A Y 
M0 Y A 0 0  TSMC18DN  L=(180E-9) W=(360E-9) AD=+1.62000000E-13 
+AS=+1.62000000E-13 PD=+1.62000000E-06 PS=+1.62000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC18DP  L=(180E-9) W=(720E-9) AD=+3.24000000E-13 
+AS=+3.24000000E-13 PD=+2.34000000E-06 PS=+2.34000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_4 
   
   
   
* FILE NAME: PROJECT_DECODER_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: DECODER.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A0 = A0
*                   A1 = A1
*                   A2 = A2
*                   NOTA0 = NOTA0
*                   NOTA1 = NOTA1
*                   NOTA2 = NOTA2
*                   W0 = W0
*                   W1 = W1
*                   W2 = W2
*                   W3 = W3
*                   W4 = W4
*                   W5 = W5
*                   W6 = W6
*                   W7 = W7
.SUBCKT DECODER_G3 A0 A1 A2 NOTA0 NOTA1 NOTA2 W0 W1 W2 W3 W4 W5 W6 W7 
XI41 A1 NOTA2 NOTA0 W2 0 VDD! NAND3_G1 
XI37 NOTA2 NOTA1 NOTA0 W0 0 VDD! NAND3_G1 
XI46 A0 NOTA2 NOTA1 W1 0 VDD! NAND3_G1 
XI48 A2 A1 A0 W7 0 VDD! NAND3_G1 
XI45 A1 A0 NOTA2 W3 0 VDD! NAND3_G1 
XI50 A2 NOTA1 NOTA0 W4 0 VDD! NAND3_G1 
XI47 A2 A0 NOTA1 W5 0 VDD! NAND3_G1 
XI49 A2 A1 NOTA0 W6 0 VDD! NAND3_G1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS DECODER_G3 
* FILE NAME: PROJECT_STAGE_1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: STAGE_1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A0 = A0
*                   A0_ = A0_
*                   A1 = A1
*                   A1_ = A1_
*                   A2 = A2
*                   A2_ = A2_
*                   CLK = CLK
*                   OUT<6> = OUT_6
*                   OUT<5> = OUT_5
*                   OUT<4> = OUT_4
*                   OUT<3> = OUT_3
*                   OUT<2> = OUT_2
*                   OUT<1> = OUT_1
*                   OUT<0> = OUT_0
*                   GND = GND
*                   VDD = VDD
.SUBCKT STAGE_1_G4 A0 A0_ A1 A1_ A2 A2_ CLK OUT_6 OUT_5 OUT_4 OUT_3 OUT_2 
+OUT_1 OUT_0 GND VDD 
XI20 CLK OUT_6 OUT_5 OUT_4 OUT_3 OUT_2 OUT_1 OUT_0 W_0 W_1 W_2 W_3 W_4 W_5 W_6 
+W_7 GND VDD MEM_8X7_G2 
XI19 A0 A1 A2 A0_ A1_ A2_ W_0 W_1 W_2 W_3 W_4 W_5 W_6 W_7 DECODER_G3 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS STAGE_1_G4 
* FILE NAME: PROJECT_NAND3_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: NAND3.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: A<2> = A_2
*                   A<1> = A_1
*                   A<0> = A_0
*                   DOUT_ = DOUT_
*                   GND = GND
*                   VDD = VDD
.SUBCKT NAND3_G1 A_2 A_1 A_0 DOUT_ GND VDD 
C3 GND A_2  45.5706E-18 M=1.0 
C4 GND A_1  36.1422E-18 M=1.0 
C5 A_0 GND  54.999E-18 M=1.0 
C6 DOUT_ VDD  76.068E-18 M=1.0 
C7 DOUT_ A_1  62.3646E-18 M=1.0 
C8 DOUT_ GND  59.4693E-18 M=1.0 
C9 DOUT_ A_0  124.7292E-18 M=1.0 
M10 DOUT_ A_0 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=449.999987495175E-9 
+AD=202.50000406976E-15 AS=121.500005152361E-15 PD=1.35000004775065E-6 
+PS=539.999973625527E-9 M=1 
M11 VDD A_1 DOUT_ VDD  TSMC18DP  L=180.000000682412E-9 W=449.999987495175E-9 
+AD=121.500005152361E-15 AS=121.500005152361E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M12 DOUT_ A_2 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=449.999987495175E-9 
+AD=121.500005152361E-15 AS=202.50000406976E-15 PD=539.999973625527E-9 
+PS=1.35000004775065E-6 M=1 
M13 DOUT_ A_0 2 GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=145.799998051317E-15 PD=1.70999999227206E-6 
+PS=360.000001364824E-9 M=1 
M14 2 A_1 1 GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M15 1 A_2 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=145.799998051317E-15 AS=364.499988352029E-15 PD=360.000001364824E-9 
+PS=1.70999999227206E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND3_G1 
* FILE NAME: PROJECT_MEM_8X7_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: MEM_8X7.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 16 12:59:16 2009.
   
* TERMINAL MAPPING: CLK = CLK
*                   OUT<6> = OUT_6
*                   OUT<5> = OUT_5
*                   OUT<4> = OUT_4
*                   OUT<3> = OUT_3
*                   OUT<2> = OUT_2
*                   OUT<1> = OUT_1
*                   OUT<0> = OUT_0
*                   W<0> = W_0
*                   W<1> = W_1
*                   W<2> = W_2
*                   W<3> = W_3
*                   W<4> = W_4
*                   W<5> = W_5
*                   W<6> = W_6
*                   W<7> = W_7
*                   GND = GND
*                   VDD = VDD
.SUBCKT MEM_8X7_G2 CLK OUT_6 OUT_5 OUT_4 OUT_3 OUT_2 OUT_1 OUT_0 W_0 W_1 W_2 
+W_3 W_4 W_5 W_6 W_7 GND VDD 
C69 GND W_6  230.9958E-18 M=1.0 
C70 GND W_5  318.9942E-18 M=1.0 
C71 GND VDD  965.23245E-18 M=1.0 
C72 GND W_4  230.9958E-18 M=1.0 
C73 GND W_3  318.9942E-18 M=1.0 
C74 CLK VDD  236.4957E-18 M=1.0 
C75 CLK GND  370.0647E-18 M=1.0 
C76 W_2 GND  230.9958E-18 M=1.0 
C77 W_1 GND  307.9944E-18 M=1.0 
C78 W_0 GND  230.9958E-18 M=1.0 
C79 W_7 GND  324.4941E-18 M=1.0 
C80 VDD OUT_2  63.8442E-18 M=1.0 
C81 OUT_1 VDD  63.8442E-18 M=1.0 
C82 W_4 14  62.3646E-18 M=1.0 
C83 OUT_0 VDD  63.8442E-18 M=1.0 
C84 GND W_6  284.2542E-18 M=1.0 
C85 GND OUT_2  125.2701E-18 M=1.0 
C86 GND W_5  370.3086E-18 M=1.0 
C87 GND VDD  2.3154021E-15 M=1.0 
C88 GND OUT_1  125.2701E-18 M=1.0 
C89 GND W_4  405.963E-18 M=1.0 
C90 GND OUT_0  125.2701E-18 M=1.0 
C91 GND W_3  492.0174E-18 M=1.0 
C92 CLK VDD  509.6133E-18 M=1.0 
C93 CLK GND  1.5018732E-15 M=1.0 
C94 W_2 GND  529.5735E-18 M=1.0 
C95 W_1 GND  685.2042E-18 M=1.0 
C96 OUT_6 VDD  63.8442E-18 M=1.0 
C97 OUT_6 GND  125.2701E-18 M=1.0 
C98 W_0 GND  668.9691E-18 M=1.0 
C99 OUT_5 VDD  63.8442E-18 M=1.0 
C100 OUT_5 GND  125.2701E-18 M=1.0 
C101 OUT_4 VDD  63.8442E-18 M=1.0 
C102 OUT_4 GND  125.2701E-18 M=1.0 
C103 W_7 49  62.3646E-18 M=1.0 
C104 W_7 48  62.3646E-18 M=1.0 
C105 W_7 45  62.3646E-18 M=1.0 
C106 W_7 44  62.3646E-18 M=1.0 
C107 W_7 42  62.3646E-18 M=1.0 
C108 W_7 GND  274.59135E-18 M=1.0 
C109 OUT_3 VDD  63.8442E-18 M=1.0 
C110 OUT_3 GND  125.2701E-18 M=1.0 
C111 W_6 50  65.0448E-18 M=1.0 
C112 W_6 48  65.0448E-18 M=1.0 
C113 W_6 45  65.0448E-18 M=1.0 
C114 W_6 44  65.0448E-18 M=1.0 
C115 W_6 43  65.0448E-18 M=1.0 
C116 W_6 42  65.0448E-18 M=1.0 
C117 W_5 52  65.0448E-18 M=1.0 
C118 W_5 51  65.0448E-18 M=1.0 
C119 W_5 41  65.0448E-18 M=1.0 
C120 W_5 40  65.0448E-18 M=1.0 
C121 W_5 39  65.0448E-18 M=1.0 
C122 W_5 38  65.0448E-18 M=1.0 
C123 W_5 W_6  110.7972E-18 M=1.0 
C124 VDD W_6  260.1792E-18 M=1.0 
C125 VDD W_5  260.1792E-18 M=1.0 
C126 W_4 55  65.0448E-18 M=1.0 
C127 W_4 54  65.0448E-18 M=1.0 
C128 W_4 37  65.0448E-18 M=1.0 
C129 W_4 18  65.0448E-18 M=1.0 
C130 W_4 17  65.0448E-18 M=1.0 
C131 W_4 14  65.0448E-18 M=1.0 
C132 W_4 W_6  110.7972E-18 M=1.0 
C133 W_4 W_5  110.7972E-18 M=1.0 
C134 W_4 VDD  1.3095432E-15 M=1.0 
C135 W_3 58  65.0448E-18 M=1.0 
C136 W_3 57  65.0448E-18 M=1.0 
C137 W_3 16  65.0448E-18 M=1.0 
C138 W_3 15  65.0448E-18 M=1.0 
C139 W_3 14  65.0448E-18 M=1.0 
C140 W_3 13  65.0448E-18 M=1.0 
C141 W_3 W_6  110.7972E-18 M=1.0 
C142 W_3 W_5  110.7972E-18 M=1.0 
C143 W_3 VDD  1.6837164E-15 M=1.0 
C144 W_3 W_4  110.7972E-18 M=1.0 
C145 GND W_6  3.6563094E-15 M=1.0 
C146 GND W_5  3.2523435E-15 M=1.0 
C147 GND W_4  3.508704E-15 M=1.0 
C148 GND W_3  1.88217E-15 M=1.0 
C149 CLK VDD  1.3826466E-15 M=1.0 
C150 CLK GND  6.75792E-15 M=1.0 
C151 W_2 61  60.31485E-18 M=1.0 
C152 W_2 60  60.31485E-18 M=1.0 
C153 W_2 12  65.0448E-18 M=1.0 
C154 W_2 11  65.0448E-18 M=1.0 
C155 W_2 10  65.0448E-18 M=1.0 
C156 W_2 9  65.0448E-18 M=1.0 
C157 W_2 W_6  110.7972E-18 M=1.0 
C158 W_2 W_5  110.7972E-18 M=1.0 
C159 W_2 VDD  874.9422E-18 M=1.0 
C160 W_2 W_4  110.7972E-18 M=1.0 
C161 W_2 W_3  110.7972E-18 M=1.0 
C162 W_2 GND  2.5909767E-15 M=1.0 
C163 W_1 64  60.31485E-18 M=1.0 
C164 W_1 63  60.31485E-18 M=1.0 
C165 W_1 8  60.31485E-18 M=1.0 
C166 W_1 7  60.31485E-18 M=1.0 
C167 W_1 6  60.31485E-18 M=1.0 
C168 W_1 5  60.31485E-18 M=1.0 
C169 W_1 W_6  110.7972E-18 M=1.0 
C170 W_1 W_5  110.7972E-18 M=1.0 
C171 W_1 VDD  874.9422E-18 M=1.0 
C172 W_1 W_4  110.7972E-18 M=1.0 
C173 W_1 W_3  110.7972E-18 M=1.0 
C174 W_1 GND  2.22498E-15 M=1.0 
C175 W_1 W_2  110.7972E-18 M=1.0 
C176 W_0 67  50.6241E-18 M=1.0 
C177 W_0 66  50.6241E-18 M=1.0 
C178 W_0 4  55.5849E-18 M=1.0 
C179 W_0 3  55.5849E-18 M=1.0 
C180 W_0 2  55.5849E-18 M=1.0 
C181 W_0 1  55.5849E-18 M=1.0 
C182 W_0 W_6  110.7972E-18 M=1.0 
C183 W_0 OUT_2  55.8603E-18 M=1.0 
C184 W_0 W_5  110.7972E-18 M=1.0 
C185 W_0 VDD  1.02615435E-15 M=1.0 
C186 W_0 OUT_1  55.62945E-18 M=1.0 
C187 W_0 W_4  110.7972E-18 M=1.0 
C188 W_0 OUT_0  55.8603E-18 M=1.0 
C189 W_0 W_3  110.7972E-18 M=1.0 
C190 W_0 GND  1.5580611E-15 M=1.0 
C191 W_0 CLK  582.5736E-18 M=1.0 
C192 W_0 W_2  110.7972E-18 M=1.0 
C193 W_0 W_1  110.7972E-18 M=1.0 
C194 OUT_5 W_0  55.62945E-18 M=1.0 
C195 OUT_4 W_0  55.8603E-18 M=1.0 
C196 W_7 48  65.0448E-18 M=1.0 
C197 W_7 47  65.0448E-18 M=1.0 
C198 W_7 46  65.0448E-18 M=1.0 
C199 W_7 45  65.0448E-18 M=1.0 
C200 W_7 44  65.0448E-18 M=1.0 
C201 W_7 42  65.0448E-18 M=1.0 
C202 W_7 W_6  110.7972E-18 M=1.0 
C203 W_7 W_5  110.7972E-18 M=1.0 
C204 W_7 VDD  260.1792E-18 M=1.0 
C205 W_7 W_4  110.7972E-18 M=1.0 
C206 W_7 W_3  110.7972E-18 M=1.0 
C207 W_7 GND  3.5733159E-15 M=1.0 
C208 W_7 W_2  110.7972E-18 M=1.0 
C209 W_7 W_1  110.7972E-18 M=1.0 
C210 W_7 W_0  110.7972E-18 M=1.0 
C211 OUT_3 W_0  55.62945E-18 M=1.0 
M212 OUT_5 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M213 OUT_3 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M214 OUT_1 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M215 VDD GND OUT_4 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M216 VDD GND OUT_2 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M217 VDD GND OUT_0 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M218 VDD GND OUT_6 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M219 VDD CLK OUT_5 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M220 VDD CLK OUT_3 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M221 VDD CLK OUT_1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M222 OUT_6 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M223 OUT_4 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M224 OUT_2 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M225 OUT_0 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M226 OUT_5 W_0 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M227 OUT_3 W_0 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M228 OUT_1 W_0 66 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M229 67 W_1 64 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M230 66 W_1 63 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M231 68 W_1 65 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M232 65 W_2 62 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M233 64 W_2 61 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M234 63 W_2 60 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M235 62 W_3 59 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M236 61 W_3 58 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M237 60 W_3 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M238 59 W_4 56 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M239 58 W_4 55 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M240 57 W_4 54 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M241 56 W_5 53 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M242 55 W_5 52 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M243 54 W_5 51 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M244 53 W_6 49 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M245 52 W_6 48 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M246 51 W_6 50 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M247 49 W_7 49 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M248 48 W_7 48 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M249 50 W_7 47 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M250 47 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M251 49 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M252 48 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M253 GND CLK 45 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M254 GND CLK 44 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M255 GND CLK 46 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M256 GND CLK 42 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M257 45 W_7 45 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M258 44 W_7 44 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M259 46 W_7 43 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M260 42 W_7 42 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M261 43 W_6 39 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M262 42 W_6 38 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M263 45 W_6 41 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M264 44 W_6 40 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M265 41 W_5 37 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M266 40 W_5 18 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M267 39 W_5 14 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M268 38 W_5 17 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M269 37 W_4 16 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M270 18 W_4 15 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M271 14 W_4 14 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M272 17 W_4 13 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M273 15 W_3 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M274 14 W_3 10 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M275 13 W_3 9 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M276 16 W_3 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M277 12 W_2 8 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M278 11 W_2 7 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M279 10 W_2 6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M280 9 W_2 5 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M281 8 W_1 4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M282 7 W_1 3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M283 6 W_1 2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M284 5 W_1 1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M285 4 W_0 OUT_6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M286 3 W_0 OUT_4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M287 2 W_0 OUT_2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M288 1 W_0 OUT_0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS MEM_8X7_G2 
   
   
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TRAN  5.00000E-11 1.50000E-08 START=  0.0000    
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
+        DELMAX = 1.00000E-10

.MEAS TRAN avg_power AVG POWER FROM=1n TO=5n
.option POST=2
.END
.END
