* # FILE NAME: /HOME/ENGR/TRUTY1/CADENCE/SIMULATION/WHOLE_CKT/HSPICES/          
* SCHEMATIC/NETLIST/WHOLE_CKT.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON DEC 8 16:24:54 2009
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: ECE482MEMORY_WHOLE_CKT_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: WHOLE_CKT.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 16:24:55 2009.
   
XI62 A0 A1 A2 CLK DFF_OUT_6 DFF_OUT_5 DFF_OUT_4 DFF_OUT_3 DFF_OUT_2 DFF_OUT_1 
+DFF_OUT_0 H_3 H_2 H_1 H_0 OUT_3 OUT_2 OUT_1 OUT_0 _DFF_OUT_6 _DFF_OUT_5 
+_DFF_OUT_4 _DFF_OUT_3 _DFF_OUT_2 _DFF_OUT_1 _DFF_OUT_0 0 VDD! PART1_G1 
C0 OUT_3 0  50E-15 M=1.0 
C3 OUT_0 0  50E-15 M=1.0 
C2 OUT_1 0  50E-15 M=1.0 
C1 OUT_2 0  50E-15 M=1.0 
VA2_GEN A2 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 6.4E-9 12.8E-9 
V1 CLK 0  PULSE 0.0 1.8 0.0 80E-12 80E-12 700E-12 1.6E-9 
VA0_GEN A0 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 1.6E-9 3.2E-9 
VA1_GEN A1 0  PULSE 1.8 0.0 -3.00000000E-10 80E-12 80E-12 3.2E-9 6.4E-9 
V0 VDD! 0  1.8 
   
   
   
   
* FILE NAME: ECE482MEMORY_PART1_EXTRACTED.S.
* SUBCIRCUIT FOR CELL: PART1.
* GENERATED FOR: HSPICES.
* GENERATED ON DEC  8 16:24:54 2009.
   
* TERMINAL MAPPING: A0 = A0
*                   A1 = A1
*                   A2 = A2
*                   CLK = CLK
*                   DFF_OUT<6> = DFF_OUT_6
*                   DFF_OUT<5> = DFF_OUT_5
*                   DFF_OUT<4> = DFF_OUT_4
*                   DFF_OUT<3> = DFF_OUT_3
*                   DFF_OUT<2> = DFF_OUT_2
*                   DFF_OUT<1> = DFF_OUT_1
*                   DFF_OUT<0> = DFF_OUT_0
*                   H<3> = H_3
*                   H<2> = H_2
*                   H<1> = H_1
*                   H<0> = H_0
*                   OUT<3> = OUT_3
*                   OUT<2> = OUT_2
*                   OUT<1> = OUT_1
*                   OUT<0> = OUT_0
*                   _DFF_OUT<6> = _DFF_OUT_6
*                   _DFF_OUT<5> = _DFF_OUT_5
*                   _DFF_OUT<4> = _DFF_OUT_4
*                   _DFF_OUT<3> = _DFF_OUT_3
*                   _DFF_OUT<2> = _DFF_OUT_2
*                   _DFF_OUT<1> = _DFF_OUT_1
*                   _DFF_OUT<0> = _DFF_OUT_0
*                   GND = GND
*                   VDD = VDD
.SUBCKT PART1_G1 A0 A1 A2 CLK DFF_OUT_6 DFF_OUT_5 DFF_OUT_4 DFF_OUT_3 
+DFF_OUT_2 DFF_OUT_1 DFF_OUT_0 H_3 H_2 H_1 H_0 OUT_3 OUT_2 OUT_1 OUT_0 
+_DFF_OUT_6 _DFF_OUT_5 _DFF_OUT_4 _DFF_OUT_3 _DFF_OUT_2 _DFF_OUT_1 _DFF_OUT_0 
+GND VDD 
C190 VDD 143  38.4992999999998E-18 M=1.0 
C191 VDD 109  280.494900000001E-18 M=1.0 
C192 VDD 102  26.7138000000001E-18 M=1.0 
C193 VDD _DFF_OUT_4  58.1418E-18 M=1.0 
C194 _DFF_OUT_2 VDD  40.0707E-18 M=1.0 
C195 GND 119  32.2137E-18 M=1.0 
C196 GND 118  32.2137E-18 M=1.0 
C197 GND 117  32.2137E-18 M=1.0 
C198 GND 116  32.2137E-18 M=1.0 
C199 GND 115  32.2137000000001E-18 M=1.0 
C200 GND 114  32.2137E-18 M=1.0 
C201 GND 113  32.2137000000001E-18 M=1.0 
C202 GND 112  318.9942E-18 M=1.0 
C203 GND _DFF_OUT_3  206.6391E-18 M=1.0 
C204 GND _DFF_OUT_2  149.283E-18 M=1.0 
C205 GND _DFF_OUT_1  206.6391E-18 M=1.0 
C206 _DFF_OUT_0 GND  206.6391E-18 M=1.0 
C207 DFF_OUT_4 GND  36.1422000000002E-18 M=1.0 
C208 _DFF_OUT_6 VDD  40.0707E-18 M=1.0 
C209 _DFF_OUT_6 GND  149.283E-18 M=1.0 
C210 112 114  62.3646E-18 M=1.0 
C211 102 111  62.3646E-18 M=1.0 
C212 95 112  62.3646E-18 M=1.0 
C213 95 111  62.3646E-18 M=1.0 
C214 67 84  62.3646E-18 M=1.0 
C215 67 76  62.3646E-18 M=1.0 
C216 67 70  62.3646E-18 M=1.0 
C217 60 70  62.3646E-18 M=1.0 
C218 28 74  62.3646E-18 M=1.0 
C219 26 84  62.3646E-18 M=1.0 
C220 16 74  62.3646E-18 M=1.0 
C221 1 81  62.3646E-18 M=1.0 
C222 1 10  62.3646E-18 M=1.0 
C223 VDD 143  46.3662000000001E-18 M=1.0 
C224 VDD 139  147.5298E-18 M=1.0 
C225 VDD 120  39.0672E-18 M=1.0 
C226 VDD 114  56.6991E-18 M=1.0 
C227 VDD 112  188.4708E-18 M=1.0 
C228 VDD 102  54.2808E-18 M=1.0 
C229 VDD 95  56.6991E-18 M=1.0 
C230 VDD 88  79.0029E-18 M=1.0 
C231 VDD 81  99.0584999999999E-18 M=1.0 
C232 VDD 10  99.0584999999998E-18 M=1.0 
C233 VDD 3  99.2619E-18 M=1.0 
C234 VDD _DFF_OUT_4  102.1419E-18 M=1.0 
C235 VDD DFF_OUT_1  54.2808E-18 M=1.0 
C236 _DFF_OUT_3 VDD  27.1404E-18 M=1.0 
C237 DFF_OUT_0 VDD  27.1404E-18 M=1.0 
C238 _DFF_OUT_2 DFF_OUT_0  62.3646E-18 M=1.0 
C239 _DFF_OUT_1 VDD  27.1404E-18 M=1.0 
C240 GND 133  448.4826E-18 M=1.0 
C241 GND 119  209.3463E-18 M=1.0 
C242 GND 118  209.3463E-18 M=1.0 
C243 GND 117  209.3463E-18 M=1.0 
C244 GND 116  209.3463E-18 M=1.0 
C245 GND 115  209.3463E-18 M=1.0 
C246 GND 114  209.3463E-18 M=1.0 
C247 GND 102  176.4513E-18 M=1.0 
C248 GND 95  195.0066E-18 M=1.0 
C249 GND 88  203.13E-18 M=1.0 
C250 GND 81  163.881E-18 M=1.0 
C251 GND 28  564.3918E-18 M=1.0 
C252 GND 10  163.881E-18 M=1.0 
C253 GND _DFF_OUT_4  267.0786E-18 M=1.0 
C254 GND _DFF_OUT_3  525.5946E-18 M=1.0 
C255 GND DFF_OUT_0  1.0597635E-15 M=1.0 
C256 GND _DFF_OUT_1  170.2845E-18 M=1.0 
C257 _DFF_OUT_0 VDD  27.1404E-18 M=1.0 
C258 _DFF_OUT_0 GND  170.2845E-18 M=1.0 
C259 _DFF_OUT_6 VDD  176.8356E-18 M=1.0 
C260 _DFF_OUT_6 DFF_OUT_4  152.442E-18 M=1.0 
C261 DFF_OUT_2 _DFF_OUT_0  62.3646E-18 M=1.0 
C262 112 114  55.3986E-18 M=1.0 
C263 102 111  104.8338E-18 M=1.0 
C264 95 111  119.3148E-18 M=1.0 
C265 95 102  297.5607E-18 M=1.0 
C266 81 109  55.3986E-18 M=1.0 
C267 67 93  65.0448E-18 M=1.0 
C268 67 84  65.0448E-18 M=1.0 
C269 67 76  65.0448E-18 M=1.0 
C270 67 70  65.0448E-18 M=1.0 
C271 60 76  65.0448E-18 M=1.0 
C272 60 70  65.0448E-18 M=1.0 
C273 28 74  65.0448E-18 M=1.0 
C274 26 93  65.0448E-18 M=1.0 
C275 26 84  65.0448E-18 M=1.0 
C276 23 28  65.0448E-18 M=1.0 
C277 16 74  64.945575E-18 M=1.0 
C278 16 21  65.0448E-18 M=1.0 
C279 10 109  55.3986E-18 M=1.0 
C280 2 74  60.31485E-18 M=1.0 
C281 2 17  60.31485E-18 M=1.0 
C282 1 81  120.3381E-18 M=1.0 
C283 1 10  120.70665E-18 M=1.0 
C284 _DFF_OUT_4 117  299.4885E-18 M=1.0 
C285 VDD 119  34.9776E-18 M=1.0 
C286 VDD 118  34.9776E-18 M=1.0 
C287 VDD 117  34.9776E-18 M=1.0 
C288 VDD 116  34.9776E-18 M=1.0 
C289 VDD 115  34.9776E-18 M=1.0 
C290 VDD 114  34.9776E-18 M=1.0 
C291 VDD 113  34.9776E-18 M=1.0 
C292 VDD 112  80.9244E-18 M=1.0 
C293 VDD 88  55.3986E-18 M=1.0 
C294 VDD 10  65.0448E-18 M=1.0 
C295 _DFF_OUT_3 116  299.4885E-18 M=1.0 
C296 _DFF_OUT_3 VDD  65.5065E-18 M=1.0 
C297 _DFF_OUT_2 115  299.4885E-18 M=1.0 
C298 _DFF_OUT_2 VDD  710.9973E-18 M=1.0 
C299 _DFF_OUT_1 114  299.4885E-18 M=1.0 
C300 _DFF_OUT_1 DFF_OUT_1  111.933E-18 M=1.0 
C301 _DFF_OUT_1 VDD  65.5065E-18 M=1.0 
C302 GND 119  48.9483E-18 M=1.0 
C303 GND 118  48.9483E-18 M=1.0 
C304 GND 117  48.9483E-18 M=1.0 
C305 GND 116  48.9483E-18 M=1.0 
C306 GND 115  48.9483E-18 M=1.0 
C307 GND 114  48.9483E-18 M=1.0 
C308 GND 113  48.9483E-18 M=1.0 
C309 GND 102  157.7223E-18 M=1.0 
C310 GND 95  107.1702E-18 M=1.0 
C311 GND 3  21.0987E-18 M=1.0 
C312 GND _DFF_OUT_4  2.7010089E-15 M=1.0 
C313 GND _DFF_OUT_3  1.3545225E-15 M=1.0 
C314 GND DFF_OUT_0  55.3986E-18 M=1.0 
C315 GND _DFF_OUT_1  537.4107E-18 M=1.0 
C316 _DFF_OUT_0 113  299.4885E-18 M=1.0 
C317 _DFF_OUT_0 _DFF_OUT_2  55.3986E-18 M=1.0 
C318 _DFF_OUT_0 GND  2.73641355E-15 M=1.0 
C319 DFF_OUT_6 _DFF_OUT_4  37.944E-18 M=1.0 
C320 DFF_OUT_4 _DFF_OUT_4  55.3986E-18 M=1.0 
C321 DFF_OUT_4 _DFF_OUT_3  55.3986E-18 M=1.0 
C322 DFF_OUT_4 _DFF_OUT_0  69.534E-18 M=1.0 
C323 _DFF_OUT_6 119  299.4885E-18 M=1.0 
C324 _DFF_OUT_6 VDD  327.7071E-18 M=1.0 
C325 _DFF_OUT_6 DFF_OUT_0  55.3986E-18 M=1.0 
C326 _DFF_OUT_6 GND  4.345002E-15 M=1.0 
C327 _DFF_OUT_6 _DFF_OUT_0  55.3986E-18 M=1.0 
C328 DFF_OUT_3 _DFF_OUT_4  110.7972E-18 M=1.0 
C329 _DFF_OUT_5 118  299.4885E-18 M=1.0 
C330 _DFF_OUT_5 DFF_OUT_5  55.3986E-18 M=1.0 
C331 DFF_OUT_2 _DFF_OUT_2  55.3986E-18 M=1.0 
C332 DFF_OUT_2 _DFF_OUT_0  69.3378E-18 M=1.0 
C333 102 112  52.3044E-18 M=1.0 
C334 95 111  37.6677E-18 M=1.0 
C335 3 109  175.510125E-18 M=1.0 
C336 3 93  104.6088E-18 M=1.0 
C337 3 88  37.6677E-18 M=1.0 
C338 3 84  104.6088E-18 M=1.0 
C339 3 81  150.907725E-18 M=1.0 
C340 3 76  104.6088E-18 M=1.0 
C341 3 70  104.6088E-18 M=1.0 
C342 3 28  104.6088E-18 M=1.0 
C343 3 16  104.6088E-18 M=1.0 
C344 3 10  163.433925E-18 M=1.0 
C345 2 3  104.6088E-18 M=1.0 
C346 1 3  104.6088E-18 M=1.0 
C347 VDD 3  388.04715E-18 M=1.0 
C348 _DFF_OUT_2 DFF_OUT_0  173.054925E-18 M=1.0 
C349 _DFF_OUT_1 _DFF_OUT_2  781.97805E-18 M=1.0 
C350 GND 139  200.52585E-18 M=1.0 
C351 GND 3  1.0969011E-15 M=1.0 
C352 GND _DFF_OUT_3  123.4143E-18 M=1.0 
C353 GND _DFF_OUT_1  1.272761775E-15 M=1.0 
C354 _DFF_OUT_0 _DFF_OUT_1  116.5779E-18 M=1.0 
C355 _DFF_OUT_0 GND  123.4143E-18 M=1.0 
C356 _DFF_OUT_6 _DFF_OUT_2  52.3044E-18 M=1.0 
C357 _DFF_OUT_6 _DFF_OUT_1  52.3044E-18 M=1.0 
C358 DFF_OUT_2 _DFF_OUT_6  52.3044E-18 M=1.0 
C359 DFF_OUT_1 133  495.25155E-18 M=1.0 
C360 _DFF_OUT_2 DFF_OUT_1  49.5477E-18 M=1.0 
C361 _DFF_OUT_6 DFF_OUT_1  49.5477E-18 M=1.0 
C362 VDD 105  26.7138E-18 M=1.0 
C363 GND 105  109.998E-18 M=1.0 
C364 GND 98  39.285E-18 M=1.0 
C365 GND 76  230.9958E-18 M=1.0 
C366 GND 70  324.4941E-18 M=1.0 
C367 GND 28  318.9942E-18 M=1.0 
C368 GND 1  230.9958E-18 M=1.0 
C369 GND VDD  958.161150000001E-18 M=1.0 
C370 112 117  62.3646E-18 M=1.0 
C371 105 111  62.3646E-18 M=1.0 
C372 98 112  62.3646E-18 M=1.0 
C373 98 111  62.3646E-18 M=1.0 
C374 73 84  62.3646E-18 M=1.0 
C375 73 76  62.3646E-18 M=1.0 
C376 68 93  62.3646E-18 M=1.0 
C377 68 84  62.3646E-18 M=1.0 
C378 68 76  62.3646E-18 M=1.0 
C379 68 70  62.3646E-18 M=1.0 
C380 1 83  62.3646E-18 M=1.0 
C381 1 82  62.3646E-18 M=1.0 
C382 VDD 117  56.6991E-18 M=1.0 
C383 VDD 111  182.6118E-18 M=1.0 
C384 VDD 109  651.0312E-18 M=1.0 
C385 VDD 105  54.2808E-18 M=1.0 
C386 VDD 98  56.6991E-18 M=1.0 
C387 VDD 89  106.7094E-18 M=1.0 
C388 VDD 83  89.3960999999999E-18 M=1.0 
C389 VDD 82  89.3961000000001E-18 M=1.0 
C390 VDD 4  72.4293E-18 M=1.0 
C391 GND 105  176.4513E-18 M=1.0 
C392 GND 98  195.0066E-18 M=1.0 
C393 GND 90  883.9386E-18 M=1.0 
C394 GND 84  442.683E-18 M=1.0 
C395 GND 83  164.9034E-18 M=1.0 
C396 GND 82  164.9034E-18 M=1.0 
C397 GND 76  349.0218E-18 M=1.0 
C398 GND 4  254.1132E-18 M=1.0 
C399 112 117  55.3986E-18 M=1.0 
C400 105 112  78.3504E-18 M=1.0 
C401 105 111  104.8338E-18 M=1.0 
C402 98 112  50.39325E-18 M=1.0 
C403 98 111  119.3148E-18 M=1.0 
C404 98 105  297.5607E-18 M=1.0 
C405 83 109  55.3986E-18 M=1.0 
C406 82 109  55.3986E-18 M=1.0 
C407 68 93  65.0448E-18 M=1.0 
C408 68 84  65.0448E-18 M=1.0 
C409 68 76  65.0448E-18 M=1.0 
C410 28 68  65.0448E-18 M=1.0 
C411 16 77  60.31485E-18 M=1.0 
C412 2 79  60.31485E-18 M=1.0 
C413 1 109  582.5736E-18 M=1.0 
C414 1 83  55.62945E-18 M=1.0 
C415 1 82  120.3381E-18 M=1.0 
C416 VDD 28  1.6542396E-15 M=1.0 
C417 VDD 5  76.4973E-18 M=1.0 
C418 GND 111  2.95639245E-15 M=1.0 
C419 GND 105  157.7223E-18 M=1.0 
C420 GND 98  107.1702E-18 M=1.0 
C421 GND 83  293.6736E-18 M=1.0 
C422 GND 82  293.6736E-18 M=1.0 
C423 GND 2  3.4484679E-15 M=1.0 
C424 105 112  52.3044E-18 M=1.0 
C425 98 111  37.6677E-18 M=1.0 
C426 5 109  156.9132E-18 M=1.0 
C427 5 90  37.6677E-18 M=1.0 
C428 5 84  104.6088E-18 M=1.0 
C429 5 83  148.216275E-18 M=1.0 
C430 5 28  104.6088E-18 M=1.0 
C431 5 16  104.6088E-18 M=1.0 
C432 4 109  156.9132E-18 M=1.0 
C433 4 93  104.6088E-18 M=1.0 
C434 4 89  37.6677E-18 M=1.0 
C435 4 82  99.2826E-18 M=1.0 
C436 4 28  138.312E-18 M=1.0 
C437 2 5  104.6088E-18 M=1.0 
C438 GND 109  326.0655E-18 M=1.0 
C439 GND 93  230.9958E-18 M=1.0 
C440 GND 84  318.9942E-18 M=1.0 
C441 GND 16  230.9958E-18 M=1.0 
C442 GND 2  307.9944E-18 M=1.0 
C443 58 76  62.3646E-18 M=1.0 
C444 57 76  62.3646E-18 M=1.0 
C445 57 70  62.3646E-18 M=1.0 
C446 25 93  62.3646E-18 M=1.0 
C447 24 93  62.3646E-18 M=1.0 
C448 19 28  62.3646E-18 M=1.0 
C449 16 19  62.3646E-18 M=1.0 
C450 16 18  62.3646E-18 M=1.0 
C451 1 13  62.3646E-18 M=1.0 
C452 1 12  62.3646E-18 M=1.0 
C453 1 11  62.3646E-18 M=1.0 
C454 VDD 13  99.0585E-18 M=1.0 
C455 VDD 12  89.3960999999999E-18 M=1.0 
C456 VDD 11  89.3961000000001E-18 M=1.0 
C457 VDD 6  81.4212E-18 M=1.0 
C458 VDD 5  74.331E-18 M=1.0 
C459 GND 93  478.3374E-18 M=1.0 
C460 GND 70  231.26985E-18 M=1.0 
C461 GND 16  601.947900000001E-18 M=1.0 
C462 GND 13  163.881E-18 M=1.0 
C463 GND 12  164.9034E-18 M=1.0 
C464 GND 11  164.9034E-18 M=1.0 
C465 GND 6  1.5927561E-15 M=1.0 
C466 GND 5  647.3034E-18 M=1.0 
C467 GND 1  741.3435E-18 M=1.0 
C468 68 70  65.0448E-18 M=1.0 
C469 63 70  65.0448E-18 M=1.0 
C470 62 70  65.0448E-18 M=1.0 
C471 61 76  65.0448E-18 M=1.0 
C472 59 84  65.0448E-18 M=1.0 
C473 58 84  65.0448E-18 M=1.0 
C474 58 76  65.0448E-18 M=1.0 
C475 57 84  65.0448E-18 M=1.0 
C476 57 76  65.0448E-18 M=1.0 
C477 57 70  65.0448E-18 M=1.0 
C478 27 93  65.0448E-18 M=1.0 
C479 25 93  65.0448E-18 M=1.0 
C480 25 28  65.0448E-18 M=1.0 
C481 24 93  65.0448E-18 M=1.0 
C482 24 28  65.0448E-18 M=1.0 
C483 19 28  65.0448E-18 M=1.0 
C484 16 22  65.0448E-18 M=1.0 
C485 16 19  65.0448E-18 M=1.0 
C486 16 18  65.0448E-18 M=1.0 
C487 13 109  55.3986E-18 M=1.0 
C488 12 109  55.3986E-18 M=1.0 
C489 11 109  55.3986E-18 M=1.0 
C490 2 20  60.31485E-18 M=1.0 
C491 2 19  60.31485E-18 M=1.0 
C492 2 18  60.31485E-18 M=1.0 
C493 1 13  64.84635E-18 M=1.0 
C494 1 12  120.70665E-18 M=1.0 
C495 1 11  120.70665E-18 M=1.0 
C496 VDD 109  1.3851225E-15 M=1.0 
C497 VDD 70  195.1344E-18 M=1.0 
C498 VDD 13  65.0448E-18 M=1.0 
C499 VDD 12  65.0448E-18 M=1.0 
C500 VDD 11  65.0448E-18 M=1.0 
C501 GND 109  5.6389419E-15 M=1.0 
C502 GND 93  4.7994795E-15 M=1.0 
C503 GND 76  4.232592E-15 M=1.0 
C504 GND 16  3.21899985E-15 M=1.0 
C505 GND 1  3.1785741E-15 M=1.0 
C506 5 93  104.6088E-18 M=1.0 
C507 5 76  104.6088E-18 M=1.0 
C508 5 70  104.6088E-18 M=1.0 
C509 5 12  161.071875E-18 M=1.0 
C510 4 84  138.312E-18 M=1.0 
C511 4 76  104.6088E-18 M=1.0 
C512 4 70  138.312E-18 M=1.0 
C513 4 16  104.6088E-18 M=1.0 
C514 4 11  113.6682E-18 M=1.0 
C515 2 4  104.6088E-18 M=1.0 
C516 1 5  104.6088E-18 M=1.0 
C517 1 4  104.6088E-18 M=1.0 
C518 VDD 5  185.822325E-18 M=1.0 
C519 VDD 4  134.736975E-18 M=1.0 
C520 GND 5  985.361175E-18 M=1.0 
C521 GND 4  973.752075E-18 M=1.0 
C522 VDD 112  271.0665E-18 M=1.0 
C523 VDD 107  26.7138E-18 M=1.0 
C524 VDD 106  26.7138E-18 M=1.0 
C525 GND 107  109.998E-18 M=1.0 
C526 GND 106  109.998E-18 M=1.0 
C527 GND 100  39.285E-18 M=1.0 
C528 GND 99  39.285E-18 M=1.0 
C529 112 119  62.3646E-18 M=1.0 
C530 112 118  62.3646E-18 M=1.0 
C531 107 111  62.3646E-18 M=1.0 
C532 106 111  62.3646E-18 M=1.0 
C533 100 112  62.3646E-18 M=1.0 
C534 100 111  62.3646E-18 M=1.0 
C535 99 112  62.3646E-18 M=1.0 
C536 99 111  62.3646E-18 M=1.0 
C537 VDD 119  56.6991E-18 M=1.0 
C538 VDD 118  56.6991E-18 M=1.0 
C539 VDD 107  54.2808E-18 M=1.0 
C540 VDD 106  54.2808E-18 M=1.0 
C541 VDD 100  56.6991E-18 M=1.0 
C542 VDD 99  56.6991E-18 M=1.0 
C543 VDD 90  81.4212E-18 M=1.0 
C544 GND 111  314.4501E-18 M=1.0 
C545 GND 107  176.4513E-18 M=1.0 
C546 GND 106  176.4513E-18 M=1.0 
C547 GND 100  195.0066E-18 M=1.0 
C548 GND 99  195.0066E-18 M=1.0 
C549 112 119  55.3986E-18 M=1.0 
C550 112 118  55.3986E-18 M=1.0 
C551 107 112  78.3504E-18 M=1.0 
C552 107 111  104.8338E-18 M=1.0 
C553 106 112  78.3504E-18 M=1.0 
C554 106 111  104.8338E-18 M=1.0 
C555 100 112  50.39325E-18 M=1.0 
C556 100 111  119.3148E-18 M=1.0 
C557 100 107  297.5607E-18 M=1.0 
C558 99 112  50.39325E-18 M=1.0 
C559 99 111  119.3148E-18 M=1.0 
C560 99 106  297.5607E-18 M=1.0 
C561 VDD 107  65.5065E-18 M=1.0 
C562 VDD 106  65.5065E-18 M=1.0 
C563 VDD 105  65.5065E-18 M=1.0 
C564 VDD 100  34.9776E-18 M=1.0 
C565 VDD 99  34.9776E-18 M=1.0 
C566 VDD 98  34.9776E-18 M=1.0 
C567 VDD 90  55.3986E-18 M=1.0 
C568 VDD 6  55.3986E-18 M=1.0 
C569 GND 107  157.7223E-18 M=1.0 
C570 GND 106  157.7223E-18 M=1.0 
C571 GND 100  107.1702E-18 M=1.0 
C572 GND 99  107.1702E-18 M=1.0 
C573 106 112  52.3044E-18 M=1.0 
C574 100 111  37.6677E-18 M=1.0 
C575 99 111  37.6677E-18 M=1.0 
C576 VDD 112  1.6100667E-15 M=1.0 
C577 VDD 111  2.24015535E-15 M=1.0 
C578 GND 112  2.2382262E-15 M=1.0 
C579 VDD 111  362.600549999999E-18 M=1.0 
C580 VDD 104  26.7138E-18 M=1.0 
C581 VDD 103  26.7138E-18 M=1.0 
C582 GND 111  288.74475E-18 M=1.0 
C583 GND 104  109.998E-18 M=1.0 
C584 GND 103  109.998E-18 M=1.0 
C585 GND 102  109.998E-18 M=1.0 
C586 GND 97  39.285E-18 M=1.0 
C587 GND 96  39.285E-18 M=1.0 
C588 GND 95  39.285E-18 M=1.0 
C589 112 116  62.3646E-18 M=1.0 
C590 112 115  62.3646E-18 M=1.0 
C591 104 111  62.3646E-18 M=1.0 
C592 103 111  62.3646E-18 M=1.0 
C593 97 112  62.3646E-18 M=1.0 
C594 97 111  62.3646E-18 M=1.0 
C595 96 112  62.3646E-18 M=1.0 
C596 96 111  62.3646E-18 M=1.0 
C597 VDD 116  56.6991E-18 M=1.0 
C598 VDD 115  56.6991E-18 M=1.0 
C599 VDD 104  54.2808E-18 M=1.0 
C600 VDD 103  54.2808E-18 M=1.0 
C601 VDD 97  56.6991E-18 M=1.0 
C602 VDD 96  56.6991E-18 M=1.0 
C603 GND 112  630.477000000001E-18 M=1.0 
C604 GND 104  176.4513E-18 M=1.0 
C605 GND 103  176.4513E-18 M=1.0 
C606 GND 97  195.0066E-18 M=1.0 
C607 GND 96  195.0066E-18 M=1.0 
C608 GND 89  460.3761E-18 M=1.0 
C609 112 116  55.3986E-18 M=1.0 
C610 112 115  55.3986E-18 M=1.0 
C611 104 112  78.3504E-18 M=1.0 
C612 104 111  104.8338E-18 M=1.0 
C613 103 112  78.3504E-18 M=1.0 
C614 103 111  104.8338E-18 M=1.0 
C615 102 112  78.3504E-18 M=1.0 
C616 97 112  50.39325E-18 M=1.0 
C617 97 111  119.3148E-18 M=1.0 
C618 97 104  297.5607E-18 M=1.0 
C619 96 112  50.39325E-18 M=1.0 
C620 96 111  119.3148E-18 M=1.0 
C621 96 103  297.5607E-18 M=1.0 
C622 95 112  50.39325E-18 M=1.0 
C623 VDD 104  65.5065E-18 M=1.0 
C624 VDD 103  65.5065E-18 M=1.0 
C625 VDD 97  34.9776E-18 M=1.0 
C626 VDD 96  34.9776E-18 M=1.0 
C627 VDD 89  55.3986E-18 M=1.0 
C628 VDD 4  73.85085E-18 M=1.0 
C629 GND 112  7.57449225000001E-15 M=1.0 
C630 GND 104  157.7223E-18 M=1.0 
C631 GND 103  157.7223E-18 M=1.0 
C632 GND 97  107.1702E-18 M=1.0 
C633 GND 96  107.1702E-18 M=1.0 
C634 104 112  52.3044E-18 M=1.0 
C635 103 112  52.3044E-18 M=1.0 
C636 97 111  37.6677E-18 M=1.0 
C637 96 111  37.6677E-18 M=1.0 
C638 VDD 110  108.426599999999E-18 M=1.0 
C639 VDD 66  53.4276E-18 M=1.0 
C640 VDD 65  139.0689E-18 M=1.0 
C641 VDD 64  53.4276000000002E-18 M=1.0 
C642 VDD 8  157.925700000001E-18 M=1.0 
C643 GND 87  204.282E-18 M=1.0 
C644 GND 72  29.8566000000003E-18 M=1.0 
C645 GND 71  29.8566000000001E-18 M=1.0 
C646 GND 65  350.422200000001E-18 M=1.0 
C647 GND 64  182.2824E-18 M=1.0 
C648 GND 8  350.422200000001E-18 M=1.0 
C649 84 86  62.3646E-18 M=1.0 
C650 76 87  124.7292E-18 M=1.0 
C651 72 110  62.3646E-18 M=1.0 
C652 71 110  62.3646000000001E-18 M=1.0 
C653 70 86  124.7292E-18 M=1.0 
C654 66 84  124.7292E-18 M=1.0 
C655 65 76  62.3646E-18 M=1.0 
C656 65 70  62.3646E-18 M=1.0 
C657 VDD 87  27.1404E-18 M=1.0 
C658 VDD 84  76.0680000000001E-18 M=1.0 
C659 VDD 76  76.0680000000001E-18 M=1.0 
C660 VDD 72  46.674E-18 M=1.0 
C661 VDD 71  46.6740000000001E-18 M=1.0 
C662 VDD 70  76.0680000000001E-18 M=1.0 
C663 VDD 66  61.8380999999999E-18 M=1.0 
C664 VDD 65  81.0251999999999E-18 M=1.0 
C665 VDD 64  54.2808000000002E-18 M=1.0 
C666 VDD 8  59.6339999999999E-18 M=1.0 
C667 VDD A1  27.1404000000001E-18 M=1.0 
C668 GND 109  1.4370291E-15 M=1.0 
C669 GND 72  205.6968E-18 M=1.0 
C670 GND 71  188.6859E-18 M=1.0 
C671 GND 66  1.4018382E-15 M=1.0 
C672 GND 65  767.791799999999E-18 M=1.0 
C673 GND 64  167.6628E-18 M=1.0 
C674 GND 8  707.1354E-18 M=1.0 
C675 GND A1  65.1743999999999E-18 M=1.0 
C676 CLK 71  62.3646000000001E-18 M=1.0 
C677 CLK 64  62.3646E-18 M=1.0 
C678 86 87  395.226E-18 M=1.0 
C679 84 93  110.7972E-18 M=1.0 
C680 84 86  146.0529E-18 M=1.0 
C681 76 93  110.7972E-18 M=1.0 
C682 76 84  110.7972E-18 M=1.0 
C683 72 110  55.3986E-18 M=1.0 
C684 71 110  75.29535E-18 M=1.0 
C685 70 93  55.3986E-18 M=1.0 
C686 70 84  55.3986E-18 M=1.0 
C687 70 76  55.3986E-18 M=1.0 
C688 66 87  55.3986E-18 M=1.0 
C689 66 86  55.3986E-18 M=1.0 
C690 66 84  55.3986E-18 M=1.0 
C691 66 76  55.3986E-18 M=1.0 
C692 66 70  55.3986E-18 M=1.0 
C693 65 87  221.5944E-18 M=1.0 
C694 65 86  221.5944E-18 M=1.0 
C695 65 76  55.93725E-18 M=1.0 
C696 65 72  345.2904E-18 M=1.0 
C697 65 70  55.93725E-18 M=1.0 
C698 65 66  55.3986E-18 M=1.0 
C699 64 110  201.6873E-18 M=1.0 
C700 64 71  342.873E-18 M=1.0 
C701 28 84  110.7972E-18 M=1.0 
C702 28 76  110.7972E-18 M=1.0 
C703 28 70  55.3986000000001E-18 M=1.0 
C704 16 84  110.7972E-18 M=1.0 
C705 16 76  110.7972E-18 M=1.0 
C706 16 70  55.3986E-18 M=1.0 
C707 16 28  110.7972E-18 M=1.0 
C708 9 87  55.3986E-18 M=1.0 
C709 9 65  55.3986E-18 M=1.0 
C710 8 87  55.3986E-18 M=1.0 
C711 8 86  55.3986E-18 M=1.0 
C712 8 84  55.3986E-18 M=1.0 
C713 8 76  55.3986E-18 M=1.0 
C714 8 70  55.3986E-18 M=1.0 
C715 8 66  221.5944E-18 M=1.0 
C716 8 65  55.3986E-18 M=1.0 
C717 8 9  311.0229E-18 M=1.0 
C718 2 84  110.7972E-18 M=1.0 
C719 2 76  110.7972E-18 M=1.0 
C720 2 70  55.3986E-18 M=1.0 
C721 2 28  110.7972E-18 M=1.0 
C722 1 84  110.7972E-18 M=1.0 
C723 1 76  110.7972E-18 M=1.0 
C724 1 70  55.3986E-18 M=1.0 
C725 1 16  110.7972E-18 M=1.0 
C726 1 2  110.7972E-18 M=1.0 
C727 VDD 93  1.3095432E-15 M=1.0 
C728 VDD 86  1.0597788E-15 M=1.0 
C729 VDD 84  260.1792E-18 M=1.0 
C730 VDD 76  260.1792E-18 M=1.0 
C731 VDD 72  34.9776E-18 M=1.0 
C732 VDD 71  34.9776E-18 M=1.0 
C733 VDD 64  65.5065E-18 M=1.0 
C734 VDD 15  34.9776E-18 M=1.0 
C735 VDD 14  34.9776E-18 M=1.0 
C736 VDD 8  445.7412E-18 M=1.0 
C737 VDD 7  65.5065E-18 M=1.0 
C738 VDD 1  1.02615435E-15 M=1.0 
C739 VDD A1  55.3986000000001E-18 M=1.0 
C740 GND 84  4.247406E-15 M=1.0 
C741 GND 72  57.4344E-18 M=1.0 
C742 GND 71  49.167E-18 M=1.0 
C743 GND 70  3.3164172E-15 M=1.0 
C744 GND 65  1.0176642E-15 M=1.0 
C745 GND 64  222.9867E-18 M=1.0 
C746 CLK 71  90.3762E-18 M=1.0 
C747 CLK 64  143.21295E-18 M=1.0 
C748 CLK VDD  1.32828435E-15 M=1.0 
C749 84 109  209.2176E-18 M=1.0 
C750 76 109  104.6088E-18 M=1.0 
C751 70 109  104.6088E-18 M=1.0 
C752 64 110  69.4476E-18 M=1.0 
C753 28 109  104.6088E-18 M=1.0 
C754 16 109  104.6088E-18 M=1.0 
C755 2 109  104.6088E-18 M=1.0 
C756 VDD 110  1.182449475E-15 M=1.0 
C757 CLK 71  52.3044000000001E-18 M=1.0 
C758 CLK 64  94.4298E-18 M=1.0 
C759 VDD 87  53.4276E-18 M=1.0 
C760 VDD 9  62.8560000000001E-18 M=1.0 
C761 GND 86  369.279000000001E-18 M=1.0 
C762 GND 66  166.5684E-18 M=1.0 
C763 GND 9  147.7116E-18 M=1.0 
C764 28 86  62.3646E-18 M=1.0 
C765 16 87  124.7292E-18 M=1.0 
C766 9 28  124.7292E-18 M=1.0 
C767 9 16  62.3646E-18 M=1.0 
C768 2 66  124.7292E-18 M=1.0 
C769 2 9  62.3646E-18 M=1.0 
C770 1 87  124.7292E-18 M=1.0 
C771 1 66  62.3646E-18 M=1.0 
C772 VDD 86  35.2638E-18 M=1.0 
C773 VDD 28  76.0680000000001E-18 M=1.0 
C774 VDD 16  76.0680000000001E-18 M=1.0 
C775 VDD 9  35.2638E-18 M=1.0 
C776 VDD 2  76.0680000000001E-18 M=1.0 
C777 VDD 1  76.0680000000001E-18 M=1.0 
C778 GND 87  1.2551877E-15 M=1.0 
C779 GND 9  771.4521E-18 M=1.0 
C780 GND 2  757.578599999999E-18 M=1.0 
C781 28 93  110.7972E-18 M=1.0 
C782 28 86  55.93725E-18 M=1.0 
C783 28 66  180.7992E-18 M=1.0 
C784 16 93  110.7972E-18 M=1.0 
C785 16 66  219.384E-18 M=1.0 
C786 9 86  55.3986E-18 M=1.0 
C787 9 66  166.1958E-18 M=1.0 
C788 9 28  55.3986E-18 M=1.0 
C789 9 16  111.33585E-18 M=1.0 
C790 2 93  110.7972E-18 M=1.0 
C791 2 66  55.3986E-18 M=1.0 
C792 2 16  110.7972E-18 M=1.0 
C793 2 9  55.3986E-18 M=1.0 
C794 1 93  110.7972E-18 M=1.0 
C795 1 66  55.3986E-18 M=1.0 
C796 1 28  110.7972E-18 M=1.0 
C797 1 9  55.3986E-18 M=1.0 
C798 VDD 65  1.0735866E-15 M=1.0 
C799 VDD 16  874.9422E-18 M=1.0 
C800 VDD 9  204.72975E-18 M=1.0 
C801 VDD 2  874.9422E-18 M=1.0 
C802 GND 87  669.15E-18 M=1.0 
C803 GND 86  922.5963E-18 M=1.0 
C804 GND 66  1.30877685E-15 M=1.0 
C805 GND 28  2.4578964E-15 M=1.0 
C806 GND 9  1.666413E-15 M=1.0 
C807 1 109  104.6088E-18 M=1.0 
C808 VDD 7  53.4276000000002E-18 M=1.0 
C809 GND 15  29.8566000000003E-18 M=1.0 
C810 GND 14  29.8566000000001E-18 M=1.0 
C811 GND 7  182.2824E-18 M=1.0 
C812 15 110  62.3646E-18 M=1.0 
C813 14 110  62.3646000000001E-18 M=1.0 
C814 VDD 15  46.674E-18 M=1.0 
C815 VDD 14  46.6740000000001E-18 M=1.0 
C816 VDD 7  54.2808000000002E-18 M=1.0 
C817 VDD A2  27.1404000000001E-18 M=1.0 
C818 GND 15  205.6968E-18 M=1.0 
C819 GND 14  188.6859E-18 M=1.0 
C820 GND 7  167.6628E-18 M=1.0 
C821 GND A2  74.6828999999998E-18 M=1.0 
C822 CLK 14  62.3646000000001E-18 M=1.0 
C823 CLK 7  62.3646E-18 M=1.0 
C824 15 110  55.3986E-18 M=1.0 
C825 14 110  75.29535E-18 M=1.0 
C826 8 15  345.2904E-18 M=1.0 
C827 7 110  201.6873E-18 M=1.0 
C828 7 14  342.873E-18 M=1.0 
C829 VDD A2  135.8802E-18 M=1.0 
C830 GND 110  2.77924995E-15 M=1.0 
C831 GND 15  57.4344E-18 M=1.0 
C832 GND 14  49.167E-18 M=1.0 
C833 GND 7  222.9867E-18 M=1.0 
C834 CLK 14  90.3762E-18 M=1.0 
C835 CLK 7  143.21295E-18 M=1.0 
C836 7 110  69.4476E-18 M=1.0 
C837 CLK 110  181.521E-18 M=1.0 
C838 CLK VDD  1.342614375E-15 M=1.0 
C839 VDD 101  26.7138000000002E-18 M=1.0 
C840 GND 101  109.998E-18 M=1.0 
C841 GND 94  39.285E-18 M=1.0 
C842 CLK GND  190.1394E-18 M=1.0 
C843 112 113  62.3646E-18 M=1.0 
C844 101 111  62.3646E-18 M=1.0 
C845 94 112  62.3646E-18 M=1.0 
C846 94 111  62.3646E-18 M=1.0 
C847 87 93  124.7292E-18 M=1.0 
C848 66 93  62.3646E-18 M=1.0 
C849 VDD 113  56.6991E-18 M=1.0 
C850 VDD 101  54.2808E-18 M=1.0 
C851 VDD 94  56.6991E-18 M=1.0 
C852 VDD 93  76.0680000000001E-18 M=1.0 
C853 GND 113  209.3463E-18 M=1.0 
C854 GND 101  176.4513E-18 M=1.0 
C855 GND 94  195.0066E-18 M=1.0 
C856 GND 3  441.8208E-18 M=1.0 
C857 CLK GND  216.0954E-18 M=1.0 
C858 112 113  55.3986E-18 M=1.0 
C859 101 112  78.3504E-18 M=1.0 
C860 101 111  104.8338E-18 M=1.0 
C861 94 112  50.39325E-18 M=1.0 
C862 94 111  119.3148E-18 M=1.0 
C863 94 101  297.5607E-18 M=1.0 
C864 3 93  233.8533E-18 M=1.0 
C865 VDD 111  2.97806175E-15 M=1.0 
C866 VDD 102  65.5065E-18 M=1.0 
C867 VDD 101  65.5065E-18 M=1.0 
C868 VDD 95  34.9776E-18 M=1.0 
C869 VDD 94  34.9776E-18 M=1.0 
C870 VDD 87  1.3209156E-15 M=1.0 
C871 VDD 66  330.2289E-18 M=1.0 
C872 VDD 3  71.2044000000001E-18 M=1.0 
C873 GND 101  157.7223E-18 M=1.0 
C874 GND 94  107.1702E-18 M=1.0 
C875 GND 81  293.6736E-18 M=1.0 
C876 GND 8  2.6106372E-15 M=1.0 
C877 GND VDD  32.1826212E-15 M=1.0 
C878 111 112  1.8995076E-15 M=1.0 
C879 101 112  52.3044E-18 M=1.0 
C880 94 111  37.6677E-18 M=1.0 
C881 93 109  209.2176E-18 M=1.0 
C882 8 109  46.2689999999999E-18 M=1.0 
C883 VDD 109  686.405475E-18 M=1.0 
C884 GND 111  1.9640457E-15 M=1.0 
C885 GND 109  2.54006685E-15 M=1.0 
C886 VDD 86  129.6405E-18 M=1.0 
C887 VDD 85  53.4276000000002E-18 M=1.0 
C888 GND 110  129.640499999998E-18 M=1.0 
C889 GND 92  29.8566000000003E-18 M=1.0 
C890 GND 91  29.8566000000001E-18 M=1.0 
C891 GND 85  182.2824E-18 M=1.0 
C892 CLK VDD  205.067699999999E-18 M=1.0 
C893 92 110  62.3646E-18 M=1.0 
C894 91 110  62.3646000000001E-18 M=1.0 
C895 VDD 110  110.7324E-18 M=1.0 
C896 VDD 108  73.3581E-18 M=1.0 
C897 VDD 92  46.674E-18 M=1.0 
C898 VDD 91  46.6740000000001E-18 M=1.0 
C899 VDD 85  54.2808000000002E-18 M=1.0 
C900 VDD A0  27.1404000000001E-18 M=1.0 
C901 GND 110  219.1122E-18 M=1.0 
C902 GND 108  144.6444E-18 M=1.0 
C903 GND 92  205.6968E-18 M=1.0 
C904 GND 91  188.6859E-18 M=1.0 
C905 GND 86  1.0601919E-15 M=1.0 
C906 GND 85  167.6628E-18 M=1.0 
C907 GND A0  76.5845999999999E-18 M=1.0 
C908 CLK 91  62.3646000000001E-18 M=1.0 
C909 CLK 85  62.3646E-18 M=1.0 
C910 CLK VDD  163.5399E-18 M=1.0 
C911 92 110  55.3986E-18 M=1.0 
C912 91 110  75.29535E-18 M=1.0 
C913 86 92  345.2904E-18 M=1.0 
C914 85 110  201.6873E-18 M=1.0 
C915 85 91  342.873E-18 M=1.0 
C916 VDD 110  65.5065E-18 M=1.0 
C917 VDD 92  34.9776E-18 M=1.0 
C918 VDD 91  34.9776E-18 M=1.0 
C919 VDD 85  65.5065E-18 M=1.0 
C920 VDD A0  55.3986000000001E-18 M=1.0 
C921 GND 92  57.4344E-18 M=1.0 
C922 GND 91  49.167E-18 M=1.0 
C923 GND 85  222.9867E-18 M=1.0 
C924 CLK 91  90.3762E-18 M=1.0 
C925 CLK 85  143.21295E-18 M=1.0 
C926 CLK GND  81.945E-18 M=1.0 
C927 85 110  69.4476E-18 M=1.0 
C928 GND 110  1.128732075E-15 M=1.0 
C929 CLK 91  52.3044000000001E-18 M=1.0 
C930 CLK 85  94.4298E-18 M=1.0 
C931 CLK GND  3.890652525E-15 M=1.0 
C932 VDD 162  40.0707E-18 M=1.0 
C933 VDD 151  220.7817E-18 M=1.0 
C934 VDD 146  38.4993E-18 M=1.0 
C935 VDD 145  38.4993E-18 M=1.0 
C936 VDD 144  38.4993E-18 M=1.0 
C937 VDD 142  51.8561999999999E-18 M=1.0 
C938 VDD 141  51.8562000000001E-18 M=1.0 
C939 VDD 140  51.8562E-18 M=1.0 
C940 VDD 139  51.8561999999999E-18 M=1.0 
C941 VDD 134  47.142E-18 M=1.0 
C942 VDD 128  58.1418E-18 M=1.0 
C943 VDD 125  21.2139000000001E-18 M=1.0 
C944 VDD DFF_OUT_1  57.945375E-18 M=1.0 
C945 GND 152  183.8538E-18 M=1.0 
C946 GND 146  58.9275E-18 M=1.0 
C947 GND 145  58.9274999999999E-18 M=1.0 
C948 GND 144  58.9275E-18 M=1.0 
C949 GND 143  58.9275000000002E-18 M=1.0 
C950 GND 142  81.7128000000001E-18 M=1.0 
C951 GND 141  81.7127999999999E-18 M=1.0 
C952 GND 140  81.7128E-18 M=1.0 
C953 GND 139  81.7127999999999E-18 M=1.0 
C954 152 158  62.3646E-18 M=1.0 
C955 150 152  62.3646E-18 M=1.0 
C956 150 151  62.3646E-18 M=1.0 
C957 149 152  62.3646E-18 M=1.0 
C958 149 151  62.3646E-18 M=1.0 
C959 148 152  62.3646E-18 M=1.0 
C960 148 151  62.3646E-18 M=1.0 
C961 147 152  62.3646E-18 M=1.0 
C962 147 151  62.3646E-18 M=1.0 
C963 131 134  62.3646E-18 M=1.0 
C964 129 142  124.7292E-18 M=1.0 
C965 128 131  62.3646E-18 M=1.0 
C966 127 142  62.3646E-18 M=1.0 
C967 125 134  62.3646E-18 M=1.0 
C968 125 131  87.1128E-18 M=1.0 
C969 DFF_OUT_1 134  62.3646E-18 M=1.0 
C970 H_2 145  124.7292E-18 M=1.0 
C971 H_2 141  124.7292E-18 M=1.0 
C972 VDD 162  27.1404E-18 M=1.0 
C973 VDD 158  56.6991E-18 M=1.0 
C974 VDD 146  46.3662E-18 M=1.0 
C975 VDD 145  46.3662E-18 M=1.0 
C976 VDD 144  46.3662E-18 M=1.0 
C977 VDD 142  147.1671E-18 M=1.0 
C978 VDD 138  39.0672E-18 M=1.0 
C979 VDD 128  48.5262E-18 M=1.0 
C980 VDD 125  151.3224E-18 M=1.0 
C981 VDD 122  27.1404E-18 M=1.0 
C982 VDD H_2  99.4158E-18 M=1.0 
C983 VDD OUT_2  47.8611E-18 M=1.0 
C984 H_1 146  124.7292E-18 M=1.0 
C985 H_1 142  124.7292E-18 M=1.0 
C986 H_1 VDD  140.2308E-18 M=1.0 
C987 _DFF_OUT_2 VDD  121.4667E-18 M=1.0 
C988 H_0 144  124.7292E-18 M=1.0 
C989 H_0 140  124.7292E-18 M=1.0 
C990 H_0 VDD  143.8803E-18 M=1.0 
C991 GND 152  264.5658E-18 M=1.0 
C992 GND 150  125.5122E-18 M=1.0 
C993 GND 149  125.5122E-18 M=1.0 
C994 GND 148  125.5122E-18 M=1.0 
C995 GND 147  125.5122E-18 M=1.0 
C996 GND 146  92.3202E-18 M=1.0 
C997 GND 145  92.3202E-18 M=1.0 
C998 GND 144  92.3202E-18 M=1.0 
C999 GND 143  92.3201999999999E-18 M=1.0 
C1000 GND 134  448.4826E-18 M=1.0 
C1001 GND 131  39.1662E-18 M=1.0 
C1002 GND 128  156.2247E-18 M=1.0 
C1003 GND 125  94.068E-18 M=1.0 
C1004 GND 122  46.1574E-18 M=1.0 
C1005 GND H_2  334.7541E-18 M=1.0 
C1006 GND H_1  268.524E-18 M=1.0 
C1007 GND H_0  308.6577E-18 M=1.0 
C1008 DFF_OUT_6 VDD  154.6749E-18 M=1.0 
C1009 DFF_OUT_6 GND  1.1417724E-15 M=1.0 
C1010 DFF_OUT_5 125  105.67395E-18 M=1.0 
C1011 DFF_OUT_5 VDD  75.3093E-18 M=1.0 
C1012 DFF_OUT_5 GND  916.66305E-18 M=1.0 
C1013 DFF_OUT_4 VDD  109.5948E-18 M=1.0 
C1014 DFF_OUT_4 GND  226.34595E-18 M=1.0 
C1015 _DFF_OUT_6 GND  261.2691E-18 M=1.0 
C1016 _DFF_OUT_5 VDD  75.0015E-18 M=1.0 
C1017 _DFF_OUT_5 GND  231.7653E-18 M=1.0 
C1018 DFF_OUT_2 VDD  124.0389E-18 M=1.0 
C1019 DFF_OUT_2 GND  706.8222E-18 M=1.0 
C1020 H_3 143  124.7292E-18 M=1.0 
C1021 H_3 139  124.7292E-18 M=1.0 
C1022 H_3 VDD  137.69145E-18 M=1.0 
C1023 H_3 GND  494.63955E-18 M=1.0 
C1024 151 154  55.3986E-18 M=1.0 
C1025 148 151  34.9776E-18 M=1.0 
C1026 142 146  59.62635E-18 M=1.0 
C1027 141 145  59.62635E-18 M=1.0 
C1028 140 144  59.62635E-18 M=1.0 
C1029 139 143  59.62635E-18 M=1.0 
C1030 128 138  74.691E-18 M=1.0 
C1031 125 131  34.9776E-18 M=1.0 
C1032 122 125  55.3986E-18 M=1.0 
C1033 _DFF_OUT_4 146  145.0206E-18 M=1.0 
C1034 _DFF_OUT_4 142  250.29945E-18 M=1.0 
C1035 _DFF_OUT_4 138  110.1303E-18 M=1.0 
C1036 _DFF_OUT_4 129  34.9776E-18 M=1.0 
C1037 _DFF_OUT_4 128  34.9776E-18 M=1.0 
C1038 _DFF_OUT_4 127  34.9776E-18 M=1.0 
C1039 H_2 145  55.3986E-18 M=1.0 
C1040 H_2 141  65.42955E-18 M=1.0 
C1041 VDD 146  250.4286E-18 M=1.0 
C1042 VDD 145  250.4286E-18 M=1.0 
C1043 VDD 144  250.4286E-18 M=1.0 
C1044 VDD 143  250.4286E-18 M=1.0 
C1045 VDD 125  130.5198E-18 M=1.0 
C1046 VDD _DFF_OUT_4  1.2171519E-15 M=1.0 
C1047 VDD H_2  135.8802E-18 M=1.0 
C1048 H_1 146  55.3986E-18 M=1.0 
C1049 H_1 142  65.42955E-18 M=1.0 
C1050 H_1 VDD  135.8802E-18 M=1.0 
C1051 _DFF_OUT_2 144  55.3986E-18 M=1.0 
C1052 _DFF_OUT_2 140  65.42955E-18 M=1.0 
C1053 H_0 144  55.3986E-18 M=1.0 
C1054 H_0 140  65.42955E-18 M=1.0 
C1055 H_0 VDD  104.5971E-18 M=1.0 
C1056 GND 165  137.0394E-18 M=1.0 
C1057 GND 151  937.6497E-18 M=1.0 
C1058 GND 146  252.9216E-18 M=1.0 
C1059 GND 145  252.9216E-18 M=1.0 
C1060 GND 144  252.9216E-18 M=1.0 
C1061 GND 143  252.9216E-18 M=1.0 
C1062 GND 142  346.2345E-18 M=1.0 
C1063 GND 141  346.2345E-18 M=1.0 
C1064 GND 140  346.2345E-18 M=1.0 
C1065 GND 139  346.2345E-18 M=1.0 
C1066 GND 125  74.1006E-18 M=1.0 
C1067 DFF_OUT_6 GND  1.4821425E-15 M=1.0 
C1068 DFF_OUT_5 134  125.3538E-18 M=1.0 
C1069 DFF_OUT_5 131  100.4841E-18 M=1.0 
C1070 DFF_OUT_5 128  65.9682E-18 M=1.0 
C1071 DFF_OUT_5 125  119.3634E-18 M=1.0 
C1072 DFF_OUT_5 122  65.9682E-18 M=1.0 
C1073 DFF_OUT_5 VDD  451.7415E-18 M=1.0 
C1074 DFF_OUT_5 GND  1.9103049E-15 M=1.0 
C1075 DFF_OUT_4 VDD  210.2778E-18 M=1.0 
C1076 DFF_OUT_4 GND  3.8796444E-15 M=1.0 
C1077 _DFF_OUT_6 143  55.3986E-18 M=1.0 
C1078 _DFF_OUT_6 139  65.42955E-18 M=1.0 
C1079 _DFF_OUT_5 145  55.3986E-18 M=1.0 
C1080 _DFF_OUT_5 141  65.42955E-18 M=1.0 
C1081 _DFF_OUT_5 VDD  1.5475599E-15 M=1.0 
C1082 _DFF_OUT_5 GND  3.4379973E-15 M=1.0 
C1083 DFF_OUT_2 DFF_OUT_1  144.1728E-18 M=1.0 
C1084 DFF_OUT_2 VDD  251.1774E-18 M=1.0 
C1085 DFF_OUT_2 GND  2.214288E-15 M=1.0 
C1086 H_3 143  55.3986E-18 M=1.0 
C1087 H_3 139  65.42955E-18 M=1.0 
C1088 H_3 VDD  135.8802E-18 M=1.0 
C1089 151 152  563.9832E-18 M=1.0 
C1090 150 151  37.6677E-18 M=1.0 
C1091 149 151  37.6677E-18 M=1.0 
C1092 148 151  37.6677E-18 M=1.0 
C1093 147 151  37.6677E-18 M=1.0 
C1094 142 146  130.1292E-18 M=1.0 
C1095 141 145  130.1292E-18 M=1.0 
C1096 140 144  130.1292E-18 M=1.0 
C1097 139 143  130.1292E-18 M=1.0 
C1098 129 142  37.6677E-18 M=1.0 
C1099 129 140  37.6677E-18 M=1.0 
C1100 128 138  114.8985E-18 M=1.0 
C1101 127 142  75.1248E-18 M=1.0 
C1102 127 128  189.8829E-18 M=1.0 
C1103 _DFF_OUT_4 129  52.3044E-18 M=1.0 
C1104 _DFF_OUT_4 128  104.6088E-18 M=1.0 
C1105 _DFF_OUT_4 127  52.3044E-18 M=1.0 
C1106 H_2 145  37.6677E-18 M=1.0 
C1107 VDD 152  384.075E-18 M=1.0 
C1108 VDD 151  1.1372994E-15 M=1.0 
C1109 VDD 146  52.3044E-18 M=1.0 
C1110 VDD 145  52.3044E-18 M=1.0 
C1111 VDD 144  52.3044E-18 M=1.0 
C1112 VDD 143  52.3044E-18 M=1.0 
C1113 VDD 142  52.3044E-18 M=1.0 
C1114 VDD 141  52.3044E-18 M=1.0 
C1115 VDD 140  52.3044E-18 M=1.0 
C1116 VDD 139  52.3044E-18 M=1.0 
C1117 H_1 146  37.6677E-18 M=1.0 
C1118 _DFF_OUT_2 129  52.3044E-18 M=1.0 
C1119 H_0 144  37.6677E-18 M=1.0 
C1120 GND 151  2.47682025E-15 M=1.0 
C1121 GND 146  278.2449E-18 M=1.0 
C1122 GND 145  278.2449E-18 M=1.0 
C1123 GND 144  278.2449E-18 M=1.0 
C1124 GND 143  278.2449E-18 M=1.0 
C1125 GND VDD  4.7622015E-15 M=1.0 
C1126 DFF_OUT_6 125  52.3044E-18 M=1.0 
C1127 DFF_OUT_6 122  155.8368E-18 M=1.0 
C1128 DFF_OUT_6 VDD  526.8573E-18 M=1.0 
C1129 DFF_OUT_5 134  33.6204E-18 M=1.0 
C1130 DFF_OUT_5 129  52.3044E-18 M=1.0 
C1131 DFF_OUT_5 128  104.6088E-18 M=1.0 
C1132 DFF_OUT_5 127  52.3044E-18 M=1.0 
C1133 DFF_OUT_5 125  211.584825E-18 M=1.0 
C1134 DFF_OUT_5 VDD  218.925675E-18 M=1.0 
C1135 DFF_OUT_5 _DFF_OUT_2  52.3044E-18 M=1.0 
C1136 DFF_OUT_5 DFF_OUT_6  52.3044E-18 M=1.0 
C1137 DFF_OUT_4 129  52.3044E-18 M=1.0 
C1138 DFF_OUT_4 DFF_OUT_5  52.3044E-18 M=1.0 
C1139 _DFF_OUT_6 128  187.6248E-18 M=1.0 
C1140 _DFF_OUT_6 DFF_OUT_5  164.53305E-18 M=1.0 
C1141 _DFF_OUT_5 125  70.614E-18 M=1.0 
C1142 _DFF_OUT_5 DFF_OUT_5  52.3044E-18 M=1.0 
C1143 DFF_OUT_2 144  173.0178E-18 M=1.0 
C1144 DFF_OUT_2 142  159.57315E-18 M=1.0 
C1145 DFF_OUT_2 140  52.3044E-18 M=1.0 
C1146 DFF_OUT_2 129  52.3044E-18 M=1.0 
C1147 DFF_OUT_2 128  52.3044E-18 M=1.0 
C1148 DFF_OUT_2 127  104.6088E-18 M=1.0 
C1149 DFF_OUT_2 _DFF_OUT_4  52.3044E-18 M=1.0 
C1150 DFF_OUT_2 VDD  577.69785E-18 M=1.0 
C1151 DFF_OUT_2 _DFF_OUT_2  104.6088E-18 M=1.0 
C1152 DFF_OUT_2 GND  1.27809585E-15 M=1.0 
C1153 DFF_OUT_2 DFF_OUT_5  52.3044E-18 M=1.0 
C1154 H_3 143  37.6677E-18 M=1.0 
C1155 VDD 135  47.142E-18 M=1.0 
C1156 VDD 129  58.1418E-18 M=1.0 
C1157 VDD 126  21.2139E-18 M=1.0 
C1158 _DFF_OUT_3 VDD  53.4276E-18 M=1.0 
C1159 GND 138  43.2135E-18 M=1.0 
C1160 GND 136  43.2135E-18 M=1.0 
C1161 GND 135  66.7845E-18 M=1.0 
C1162 GND 134  66.7845000000001E-18 M=1.0 
C1163 GND 132  58.9275E-18 M=1.0 
C1164 GND 131  58.9275000000001E-18 M=1.0 
C1165 GND 129  174.4254E-18 M=1.0 
C1166 GND 128  136.7118E-18 M=1.0 
C1167 GND 127  127.2834E-18 M=1.0 
C1168 GND 126  27.4995E-18 M=1.0 
C1169 GND 125  27.4995E-18 M=1.0 
C1170 DFF_OUT_5 VDD  155.96145E-18 M=1.0 
C1171 DFF_OUT_5 GND  73.46295E-18 M=1.0 
C1172 DFF_OUT_3 VDD  65.2131E-18 M=1.0 
C1173 DFF_OUT_3 GND  52.6419E-18 M=1.0 
C1174 _DFF_OUT_5 VDD  77.7843000000001E-18 M=1.0 
C1175 _DFF_OUT_5 GND  252.9954E-18 M=1.0 
C1176 132 135  62.3646E-18 M=1.0 
C1177 129 132  62.3646E-18 M=1.0 
C1178 128 140  124.7292E-18 M=1.0 
C1179 127 140  62.3646E-18 M=1.0 
C1180 126 135  62.3646E-18 M=1.0 
C1181 126 132  87.1128E-18 M=1.0 
C1182 VDD 140  147.1671E-18 M=1.0 
C1183 VDD 136  39.0672E-18 M=1.0 
C1184 VDD 135  69.4944E-18 M=1.0 
C1185 VDD 129  38.99025E-18 M=1.0 
C1186 VDD 126  151.3224E-18 M=1.0 
C1187 VDD 123  27.1404E-18 M=1.0 
C1188 _DFF_OUT_3 135  62.3646E-18 M=1.0 
C1189 GND 142  151.0308E-18 M=1.0 
C1190 GND 140  151.0308E-18 M=1.0 
C1191 GND 138  75.6612E-18 M=1.0 
C1192 GND 136  156.58695E-18 M=1.0 
C1193 GND 135  448.4826E-18 M=1.0 
C1194 GND 132  39.1662E-18 M=1.0 
C1195 GND 129  185.83875E-18 M=1.0 
C1196 GND 127  130.167E-18 M=1.0 
C1197 GND 126  94.068E-18 M=1.0 
C1198 GND 123  46.1574E-18 M=1.0 
C1199 DFF_OUT_5 126  105.67395E-18 M=1.0 
C1200 DFF_OUT_4 _DFF_OUT_3  62.3646E-18 M=1.0 
C1201 DFF_OUT_3 135  62.3646E-18 M=1.0 
C1202 DFF_OUT_3 _DFF_OUT_4  62.3646E-18 M=1.0 
C1203 DFF_OUT_3 VDD  32.6421E-18 M=1.0 
C1204 DFF_OUT_3 GND  371.5074E-18 M=1.0 
C1205 _DFF_OUT_5 126  62.3646E-18 M=1.0 
C1206 _DFF_OUT_5 DFF_OUT_6  124.7292E-18 M=1.0 
C1207 129 136  20.7792E-18 M=1.0 
C1208 129 135  90.3762E-18 M=1.0 
C1209 129 132  100.40715E-18 M=1.0 
C1210 128 140  166.1958E-18 M=1.0 
C1211 128 136  34.9776E-18 M=1.0 
C1212 128 134  90.3762E-18 M=1.0 
C1213 128 131  100.4841E-18 M=1.0 
C1214 128 129  20.7792E-18 M=1.0 
C1215 127 129  20.7792E-18 M=1.0 
C1216 127 128  34.9776E-18 M=1.0 
C1217 126 132  34.9776E-18 M=1.0 
C1218 126 129  120.82815E-18 M=1.0 
C1219 125 128  120.9051E-18 M=1.0 
C1220 123 126  55.3986E-18 M=1.0 
C1221 _DFF_OUT_4 134  113.2758E-18 M=1.0 
C1222 VDD 128  488.2302E-18 M=1.0 
C1223 VDD 126  130.5198E-18 M=1.0 
C1224 _DFF_OUT_3 _DFF_OUT_4  55.3986E-18 M=1.0 
C1225 GND 129  1.2261537E-15 M=1.0 
C1226 GND 128  852.8643E-18 M=1.0 
C1227 GND 126  74.1006E-18 M=1.0 
C1228 GND _DFF_OUT_2  4.2521103E-15 M=1.0 
C1229 DFF_OUT_5 _DFF_OUT_4  55.3986E-18 M=1.0 
C1230 DFF_OUT_5 _DFF_OUT_3  55.3986E-18 M=1.0 
C1231 DFF_OUT_4 142  60.46875E-18 M=1.0 
C1232 DFF_OUT_4 138  34.9776E-18 M=1.0 
C1233 DFF_OUT_4 135  60.165E-18 M=1.0 
C1234 DFF_OUT_4 129  34.9776E-18 M=1.0 
C1235 DFF_OUT_4 127  34.9776E-18 M=1.0 
C1236 _DFF_OUT_6 126  89.48835E-18 M=1.0 
C1237 _DFF_OUT_6 DFF_OUT_6  171.26595E-18 M=1.0 
C1238 _DFF_OUT_6 DFF_OUT_5  133.3746E-18 M=1.0 
C1239 DFF_OUT_3 135  55.3986E-18 M=1.0 
C1240 DFF_OUT_3 134  299.3148E-18 M=1.0 
C1241 DFF_OUT_3 _DFF_OUT_3  187.5924E-18 M=1.0 
C1242 DFF_OUT_3 GND  1.0568331E-15 M=1.0 
C1243 DFF_OUT_3 DFF_OUT_5  55.3986E-18 M=1.0 
C1244 DFF_OUT_3 DFF_OUT_4  258.642E-18 M=1.0 
C1245 _DFF_OUT_5 DFF_OUT_6  131.2866E-18 M=1.0 
C1246 127 140  75.6513E-18 M=1.0 
C1247 VDD _DFF_OUT_4  189.830025E-18 M=1.0 
C1248 _DFF_OUT_3 VDD  52.3044E-18 M=1.0 
C1249 _DFF_OUT_2 128  104.6088E-18 M=1.0 
C1250 _DFF_OUT_2 _DFF_OUT_4  52.3044E-18 M=1.0 
C1251 GND 140  44.1036E-18 M=1.0 
C1252 GND 138  37.6677E-18 M=1.0 
C1253 GND 136  192.4263E-18 M=1.0 
C1254 GND 129  1.780714575E-15 M=1.0 
C1255 DFF_OUT_6 _DFF_OUT_3  52.3044E-18 M=1.0 
C1256 DFF_OUT_6 GND  639.31725E-18 M=1.0 
C1257 DFF_OUT_5 _DFF_OUT_4  104.6088E-18 M=1.0 
C1258 DFF_OUT_5 _DFF_OUT_3  52.3044E-18 M=1.0 
C1259 DFF_OUT_5 GND  392.5071E-18 M=1.0 
C1260 DFF_OUT_4 128  153.4293E-18 M=1.0 
C1261 DFF_OUT_4 127  104.6088E-18 M=1.0 
C1262 DFF_OUT_4 _DFF_OUT_4  156.9132E-18 M=1.0 
C1263 DFF_OUT_4 VDD  312.459525E-18 M=1.0 
C1264 DFF_OUT_4 _DFF_OUT_2  156.9132E-18 M=1.0 
C1265 DFF_OUT_4 GND  1.3126095E-15 M=1.0 
C1266 _DFF_OUT_6 126  150.1443E-18 M=1.0 
C1267 _DFF_OUT_6 VDD  368.2359E-18 M=1.0 
C1268 _DFF_OUT_6 _DFF_OUT_3  52.3044E-18 M=1.0 
C1269 DFF_OUT_3 VDD  52.3044E-18 M=1.0 
C1270 DFF_OUT_3 DFF_OUT_6  52.3044E-18 M=1.0 
C1271 DFF_OUT_3 DFF_OUT_5  52.3044E-18 M=1.0 
C1272 DFF_OUT_3 DFF_OUT_4  227.9799E-18 M=1.0 
C1273 DFF_OUT_3 _DFF_OUT_6  52.3044E-18 M=1.0 
C1274 _DFF_OUT_5 _DFF_OUT_4  52.3044E-18 M=1.0 
C1275 _DFF_OUT_5 _DFF_OUT_3  52.3044E-18 M=1.0 
C1276 _DFF_OUT_5 _DFF_OUT_6  140.1714E-18 M=1.0 
C1277 _DFF_OUT_5 DFF_OUT_3  52.3044E-18 M=1.0 
C1278 VDD 133  47.1419999999999E-18 M=1.0 
C1279 VDD 127  58.1418E-18 M=1.0 
C1280 VDD 124  21.2139E-18 M=1.0 
C1281 DFF_OUT_0 VDD  57.9453750000001E-18 M=1.0 
C1282 _DFF_OUT_1 VDD  53.4276000000001E-18 M=1.0 
C1283 GND 137  43.2135E-18 M=1.0 
C1284 GND 133  66.7845000000001E-18 M=1.0 
C1285 GND 130  58.9275000000004E-18 M=1.0 
C1286 GND 124  27.4995000000001E-18 M=1.0 
C1287 GND _DFF_OUT_4  201.9249E-18 M=1.0 
C1288 GND DFF_OUT_1  59.9096249999999E-18 M=1.0 
C1289 GND DFF_OUT_0  59.909625E-18 M=1.0 
C1290 _DFF_OUT_0 VDD  53.4276000000002E-18 M=1.0 
C1291 DFF_OUT_4 VDD  78.5699999999998E-18 M=1.0 
C1292 130 133  62.3646E-18 M=1.0 
C1293 129 141  124.7292E-18 M=1.0 
C1294 129 139  124.7292E-18 M=1.0 
C1295 128 141  62.3646E-18 M=1.0 
C1296 128 139  62.3646E-18 M=1.0 
C1297 127 130  62.3646E-18 M=1.0 
C1298 124 133  62.3646E-18 M=1.0 
C1299 124 130  87.1128E-18 M=1.0 
C1300 _DFF_OUT_4 124  62.3646E-18 M=1.0 
C1301 VDD 141  147.1671E-18 M=1.0 
C1302 VDD 137  39.0672E-18 M=1.0 
C1303 VDD 134  69.4944E-18 M=1.0 
C1304 VDD 133  69.4944E-18 M=1.0 
C1305 VDD 127  41.6889E-18 M=1.0 
C1306 VDD 124  151.3224E-18 M=1.0 
C1307 VDD 121  27.1404E-18 M=1.0 
C1308 DFF_OUT_0 133  62.3646E-18 M=1.0 
C1309 _DFF_OUT_2 DFF_OUT_1  62.3646E-18 M=1.0 
C1310 _DFF_OUT_1 134  62.3646E-18 M=1.0 
C1311 GND 141  151.0308E-18 M=1.0 
C1312 GND 139  152.262E-18 M=1.0 
C1313 GND 137  75.6612E-18 M=1.0 
C1314 GND 130  39.1662E-18 M=1.0 
C1315 GND 124  94.068E-18 M=1.0 
C1316 GND 121  46.1574E-18 M=1.0 
C1317 GND DFF_OUT_1  467.829000000001E-18 M=1.0 
C1318 GND _DFF_OUT_2  432.1692E-18 M=1.0 
C1319 _DFF_OUT_0 133  62.3646E-18 M=1.0 
C1320 DFF_OUT_6 _DFF_OUT_4  62.3646E-18 M=1.0 
C1321 DFF_OUT_4 124  105.67395E-18 M=1.0 
C1322 _DFF_OUT_6 DFF_OUT_5  304.884E-18 M=1.0 
C1323 _DFF_OUT_5 125  62.3646E-18 M=1.0 
C1324 DFF_OUT_2 _DFF_OUT_1  62.3646E-18 M=1.0 
C1325 128 137  114.4917E-18 M=1.0 
C1326 127 133  90.3762E-18 M=1.0 
C1327 127 130  100.40715E-18 M=1.0 
C1328 124 130  34.9776E-18 M=1.0 
C1329 124 127  120.82815E-18 M=1.0 
C1330 121 124  55.3986E-18 M=1.0 
C1331 DFF_OUT_1 134  73.8648E-18 M=1.0 
C1332 VDD 133  55.3986E-18 M=1.0 
C1333 VDD 127  797.38335E-18 M=1.0 
C1334 VDD 124  130.5198E-18 M=1.0 
C1335 VDD DFF_OUT_1  47.74545E-18 M=1.0 
C1336 _DFF_OUT_2 DFF_OUT_1  55.3986E-18 M=1.0 
C1337 GND 127  576.7623E-18 M=1.0 
C1338 GND 124  74.1006E-18 M=1.0 
C1339 GND DFF_OUT_1  43.10865E-18 M=1.0 
C1340 _DFF_OUT_0 124  133.87995E-18 M=1.0 
C1341 _DFF_OUT_0 _DFF_OUT_4  59.436E-18 M=1.0 
C1342 _DFF_OUT_0 VDD  192.4776E-18 M=1.0 
C1343 DFF_OUT_6 133  125.3538E-18 M=1.0 
C1344 DFF_OUT_6 130  100.4841E-18 M=1.0 
C1345 DFF_OUT_6 127  65.9682E-18 M=1.0 
C1346 DFF_OUT_6 124  65.5065E-18 M=1.0 
C1347 DFF_OUT_6 121  85.6575E-18 M=1.0 
C1348 DFF_OUT_6 VDD  245.3391E-18 M=1.0 
C1349 DFF_OUT_6 _DFF_OUT_0  134.75475E-18 M=1.0 
C1350 DFF_OUT_4 133  380.68425E-18 M=1.0 
C1351 _DFF_OUT_6 125  65.2635E-18 M=1.0 
C1352 _DFF_OUT_6 124  65.2635E-18 M=1.0 
C1353 _DFF_OUT_6 _DFF_OUT_4  49.176E-18 M=1.0 
C1354 _DFF_OUT_6 DFF_OUT_4  49.1985E-18 M=1.0 
C1355 _DFF_OUT_5 137  75.1527E-18 M=1.0 
C1356 _DFF_OUT_5 127  34.9776E-18 M=1.0 
C1357 _DFF_OUT_5 _DFF_OUT_6  98.352E-18 M=1.0 
C1358 DFF_OUT_2 134  94.2021E-18 M=1.0 
C1359 DFF_OUT_2 133  60.165E-18 M=1.0 
C1360 DFF_OUT_2 DFF_OUT_0  49.176E-18 M=1.0 
C1361 129 141  148.71645E-18 M=1.0 
C1362 129 137  51.0561E-18 M=1.0 
C1363 128 137  111.78585E-18 M=1.0 
C1364 128 129  25.6374E-18 M=1.0 
C1365 VDD 129  640.033875E-18 M=1.0 
C1366 VDD 128  235.9845E-18 M=1.0 
C1367 VDD 127  219.86595E-18 M=1.0 
C1368 _DFF_OUT_2 127  104.6088E-18 M=1.0 
C1369 _DFF_OUT_2 DFF_OUT_1  194.900625E-18 M=1.0 
C1370 _DFF_OUT_2 VDD  122.9121E-18 M=1.0 
C1371 _DFF_OUT_1 133  93.7305E-18 M=1.0 
C1372 _DFF_OUT_1 130  141.3855E-18 M=1.0 
C1373 _DFF_OUT_1 127  52.3044E-18 M=1.0 
C1374 _DFF_OUT_1 VDD  307.445175E-18 M=1.0 
C1375 GND 137  37.6677E-18 M=1.0 
C1376 GND 128  1.1781747E-15 M=1.0 
C1377 GND 127  1.218818925E-15 M=1.0 
C1378 GND _DFF_OUT_4  2.242333575E-15 M=1.0 
C1379 GND _DFF_OUT_2  1.52013015E-15 M=1.0 
C1380 _DFF_OUT_0 _DFF_OUT_4  52.3044E-18 M=1.0 
C1381 DFF_OUT_6 129  52.3044E-18 M=1.0 
C1382 DFF_OUT_6 128  52.3044E-18 M=1.0 
C1383 DFF_OUT_6 127  52.3044E-18 M=1.0 
C1384 DFF_OUT_6 124  52.3044E-18 M=1.0 
C1385 DFF_OUT_6 121  141.435E-18 M=1.0 
C1386 DFF_OUT_6 _DFF_OUT_4  57.4173E-18 M=1.0 
C1387 DFF_OUT_6 _DFF_OUT_2  52.3044E-18 M=1.0 
C1388 DFF_OUT_6 _DFF_OUT_1  52.3044E-18 M=1.0 
C1389 DFF_OUT_6 _DFF_OUT_0  119.8719E-18 M=1.0 
C1390 DFF_OUT_4 124  231.738075E-18 M=1.0 
C1391 DFF_OUT_4 DFF_OUT_1  51.138E-18 M=1.0 
C1392 DFF_OUT_4 _DFF_OUT_1  52.3044E-18 M=1.0 
C1393 DFF_OUT_4 DFF_OUT_6  104.6088E-18 M=1.0 
C1394 _DFF_OUT_6 127  187.6248E-18 M=1.0 
C1395 _DFF_OUT_6 125  252.9882E-18 M=1.0 
C1396 _DFF_OUT_6 124  181.39725E-18 M=1.0 
C1397 _DFF_OUT_6 _DFF_OUT_4  86.9805E-18 M=1.0 
C1398 _DFF_OUT_6 GND  694.307475E-18 M=1.0 
C1399 _DFF_OUT_6 _DFF_OUT_0  128.8809E-18 M=1.0 
C1400 _DFF_OUT_6 DFF_OUT_6  52.3044E-18 M=1.0 
C1401 _DFF_OUT_6 DFF_OUT_4  136.78245E-18 M=1.0 
C1402 _DFF_OUT_5 129  52.3044E-18 M=1.0 
C1403 _DFF_OUT_5 128  132.0732E-18 M=1.0 
C1404 _DFF_OUT_5 127  52.3044E-18 M=1.0 
C1405 _DFF_OUT_5 VDD  530.63775E-18 M=1.0 
C1406 _DFF_OUT_5 _DFF_OUT_2  52.3044E-18 M=1.0 
C1407 _DFF_OUT_5 _DFF_OUT_1  52.3044E-18 M=1.0 
C1408 _DFF_OUT_5 GND  817.0281E-18 M=1.0 
C1409 _DFF_OUT_5 DFF_OUT_6  114.8346E-18 M=1.0 
C1410 _DFF_OUT_5 DFF_OUT_4  52.3044E-18 M=1.0 
C1411 DFF_OUT_2 133  56.3436E-18 M=1.0 
C1412 DFF_OUT_2 DFF_OUT_0  51.110775E-18 M=1.0 
C1413 DFF_OUT_2 _DFF_OUT_1  180.868725E-18 M=1.0 
C1414 DFF_OUT_2 DFF_OUT_6  52.3044E-18 M=1.0 
C1415 DFF_OUT_2 DFF_OUT_4  156.9132E-18 M=1.0 
C1416 DFF_OUT_2 _DFF_OUT_5  52.3044E-18 M=1.0 
C1417 DFF_OUT_1 134  87.12585E-18 M=1.0 
C1418 DFF_OUT_1 127  49.5477E-18 M=1.0 
C1419 VDD DFF_OUT_1  179.4771E-18 M=1.0 
C1420 GND DFF_OUT_1  823.8654E-18 M=1.0 
C1421 _DFF_OUT_0 DFF_OUT_1  75.5973E-18 M=1.0 
C1422 DFF_OUT_6 DFF_OUT_1  49.5477E-18 M=1.0 
C1423 DFF_OUT_4 DFF_OUT_1  49.5477E-18 M=1.0 
C1424 _DFF_OUT_5 DFF_OUT_1  49.5477E-18 M=1.0 
C1425 VDD 164  40.0707E-18 M=1.0 
C1426 VDD 163  40.0707E-18 M=1.0 
C1427 GND 164  148.4973E-18 M=1.0 
C1428 GND 163  148.4973E-18 M=1.0 
C1429 GND 160  38.4993E-18 M=1.0 
C1430 GND 159  38.4993E-18 M=1.0 
C1431 GND 151  173.6397E-18 M=1.0 
C1432 GND 150  38.4993E-18 M=1.0 
C1433 GND 149  38.4993E-18 M=1.0 
C1434 152 160  62.3646E-18 M=1.0 
C1435 152 159  62.3646E-18 M=1.0 
C1436 151 156  62.3646E-18 M=1.0 
C1437 151 155  62.3646E-18 M=1.0 
C1438 VDD 164  27.1404E-18 M=1.0 
C1439 VDD 163  27.1404E-18 M=1.0 
C1440 VDD 160  56.6991E-18 M=1.0 
C1441 VDD 159  56.6991E-18 M=1.0 
C1442 VDD 156  54.2808E-18 M=1.0 
C1443 VDD 155  54.2808E-18 M=1.0 
C1444 VDD 151  168.6348E-18 M=1.0 
C1445 OUT_1 VDD  47.8611E-18 M=1.0 
C1446 OUT_0 VDD  47.8611E-18 M=1.0 
C1447 GND 164  162.0072E-18 M=1.0 
C1448 GND 163  162.0072E-18 M=1.0 
C1449 GND 160  226.4616E-18 M=1.0 
C1450 GND 159  226.4616E-18 M=1.0 
C1451 GND 156  120.8403E-18 M=1.0 
C1452 GND 155  120.8403E-18 M=1.0 
C1453 GND 151  189.7794E-18 M=1.0 
C1454 GND VDD  5.88871935E-15 M=1.0 
C1455 GND OUT_1  98.3826E-18 M=1.0 
C1456 GND OUT_0  98.3826E-18 M=1.0 
C1457 160 164  306.8514E-18 M=1.0 
C1458 159 163  306.8514E-18 M=1.0 
C1459 152 160  120.9051E-18 M=1.0 
C1460 152 159  120.9051E-18 M=1.0 
C1461 152 156  230.1192E-18 M=1.0 
C1462 152 155  230.1192E-18 M=1.0 
C1463 151 156  55.3986E-18 M=1.0 
C1464 151 155  55.3986E-18 M=1.0 
C1465 151 152  139.9104E-18 M=1.0 
C1466 150 152  49.176E-18 M=1.0 
C1467 150 151  34.9776E-18 M=1.0 
C1468 149 152  49.176E-18 M=1.0 
C1469 149 151  34.9776E-18 M=1.0 
C1470 OUT_1 163  55.3986E-18 M=1.0 
C1471 OUT_0 164  55.3986E-18 M=1.0 
C1472 GND 164  559.068525E-18 M=1.0 
C1473 GND 163  559.068525E-18 M=1.0 
C1474 GND 160  113.0463E-18 M=1.0 
C1475 GND 159  113.0463E-18 M=1.0 
C1476 GND 152  1.9858005E-15 M=1.0 
C1477 150 152  212.5242E-18 M=1.0 
C1478 149 152  212.5242E-18 M=1.0 
C1479 VDD 161  40.0707E-18 M=1.0 
C1480 VDD 152  133.569E-18 M=1.0 
C1481 GND 162  148.4973E-18 M=1.0 
C1482 GND 161  148.4973E-18 M=1.0 
C1483 GND 158  38.4993E-18 M=1.0 
C1484 GND 157  38.4993000000001E-18 M=1.0 
C1485 GND 148  38.4993E-18 M=1.0 
C1486 GND 147  38.4993000000001E-18 M=1.0 
C1487 152 157  62.3646E-18 M=1.0 
C1488 151 154  62.3646E-18 M=1.0 
C1489 151 153  62.3646E-18 M=1.0 
C1490 VDD 161  27.1404E-18 M=1.0 
C1491 VDD 157  56.6991E-18 M=1.0 
C1492 VDD 154  54.2808E-18 M=1.0 
C1493 VDD 153  54.2808E-18 M=1.0 
C1494 VDD 152  67.0428E-18 M=1.0 
C1495 GND 162  162.0072E-18 M=1.0 
C1496 GND 161  162.0072E-18 M=1.0 
C1497 GND 158  226.4616E-18 M=1.0 
C1498 GND 157  226.4616E-18 M=1.0 
C1499 GND 154  120.8403E-18 M=1.0 
C1500 GND 153  120.8403E-18 M=1.0 
C1501 GND OUT_2  98.3826E-18 M=1.0 
C1502 OUT_3 VDD  47.8611E-18 M=1.0 
C1503 OUT_3 GND  98.3826E-18 M=1.0 
C1504 158 162  306.8514E-18 M=1.0 
C1505 157 161  306.8514E-18 M=1.0 
C1506 152 158  120.9051E-18 M=1.0 
C1507 152 157  120.9051E-18 M=1.0 
C1508 152 154  230.1192E-18 M=1.0 
C1509 152 153  230.1192E-18 M=1.0 
C1510 151 153  55.3986E-18 M=1.0 
C1511 148 152  49.176E-18 M=1.0 
C1512 147 152  49.176E-18 M=1.0 
C1513 147 151  34.9776E-18 M=1.0 
C1514 OUT_2 162  55.3986E-18 M=1.0 
C1515 GND 162  559.068525E-18 M=1.0 
C1516 GND 161  559.068525E-18 M=1.0 
C1517 GND 158  113.0463E-18 M=1.0 
C1518 GND 157  113.0463E-18 M=1.0 
C1519 OUT_3 161  55.3986E-18 M=1.0 
C1520 148 152  212.5242E-18 M=1.0 
C1521 147 152  212.5242E-18 M=1.0 
C1522 GND 152  2.432469375E-15 M=1.0 
C1523 GND 120  38.4993000000001E-18 M=1.0 
C1524 GND 120  1.10029275E-15 M=1.0 
C1525 VDD 152  60.46875E-18 M=1.0 
C1526 VDD 151  1.39076235E-15 M=1.0 
C1527 VDD 120  90.3762E-18 M=1.0 
C1528 GND 120  261.0576E-18 M=1.0 
C1529 _DFF_OUT_0 DFF_OUT_1  55.3986E-18 M=1.0 
C1530 _DFF_OUT_0 DFF_OUT_0  110.7972E-18 M=1.0 
M1531 83 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1532 82 GND VDD VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1533 VDD GND 10 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1534 VDD GND 13 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1535 VDD GND 12 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1536 VDD GND 11 VDD  TSMC18DP  L=1.35000004775065E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1537 81 GND VDD VDD  TSMC18DP  L=1.17000001864653E-6 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1538 87 86 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1539 66 65 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1540 9 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1541 93 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1542 VDD 66 93 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1543 93 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1544 84 66 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1545 VDD 86 84 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1546 84 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1547 76 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1548 VDD 65 76 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1549 76 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1550 70 86 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1551 VDD 65 70 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1552 70 8 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1553 28 9 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1554 VDD 86 28 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1555 28 65 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1556 16 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1557 VDD 9 16 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1558 16 65 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1559 2 66 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1560 VDD 9 2 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1561 2 86 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1562 1 87 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=283.500002987158E-15 AS=170.1000045028E-15 PD=1.52999996316794E-6 
+PS=539.999973625527E-9 M=1 
M1563 VDD 66 1 VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=170.1000045028E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1564 1 9 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=629.999988177588E-9 
+AD=170.1000045028E-15 AS=283.500002987158E-15 PD=539.999973625527E-9 
+PS=1.52999996316794E-6 M=1 
M1565 91 CLK A0 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1566 71 CLK A1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1567 14 CLK A2 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1568 85 91 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1569 86 92 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1570 65 72 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1571 64 71 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1572 8 15 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1573 7 14 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=3.24000006912684E-6 
+AD=1.45799995340812E-12 AS=1.45799995340812E-12 PD=4.13999987358693E-6 
+PS=4.13999987358693E-6 M=1 
M1574 92 110 85 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1575 72 110 64 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1576 15 110 7 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1577 92 86 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1578 91 85 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1579 72 65 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1580 71 64 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1581 15 8 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1582 14 7 VDD VDD  TSMC18DP  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1583 109 108 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1584 108 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1585 112 111 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1586 111 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1587 110 CLK VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1588 _DFF_OUT_6 119 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1589 _DFF_OUT_5 118 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1590 _DFF_OUT_4 117 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1591 _DFF_OUT_3 116 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1592 _DFF_OUT_2 115 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1593 _DFF_OUT_1 114 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1594 _DFF_OUT_0 113 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=2.70000009550131E-6 AD=1.2149999973135E-12 AS=1.2149999973135E-12 
+PD=3.5999998999614E-6 PS=3.5999998999614E-6 M=1 
M1595 DFF_OUT_3 _DFF_OUT_3 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1596 DFF_OUT_2 _DFF_OUT_2 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1597 DFF_OUT_1 _DFF_OUT_1 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1598 DFF_OUT_0 _DFF_OUT_0 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1599 DFF_OUT_6 _DFF_OUT_6 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1600 DFF_OUT_5 _DFF_OUT_5 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1601 DFF_OUT_4 _DFF_OUT_4 VDD VDD  TSMC18DP  L=180.000000682412E-9 
+W=1.62000003456342E-6 AD=728.999976704059E-15 AS=728.999976704059E-15 
+PD=2.51999995271035E-6 PS=2.51999995271035E-6 M=1 
M1602 107 100 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1603 106 99 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1604 105 98 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1605 104 97 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1606 103 96 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1607 102 95 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1608 101 94 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1609 146 142 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1610 145 141 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1611 144 140 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1612 143 139 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1613 142 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1614 141 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1615 140 128 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1616 VDD 127 142 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1617 VDD 128 141 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1618 VDD 127 140 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1619 142 138 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1620 141 137 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1621 139 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1622 140 136 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1623 VDD 128 139 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1624 138 128 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1625 137 127 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1626 139 127 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1627 136 129 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1628 _DFF_OUT_4 _DFF_OUT_3 135 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1629 _DFF_OUT_2 _DFF_OUT_1 134 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1630 _DFF_OUT_2 _DFF_OUT_0 133 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1631 135 DFF_OUT_3 DFF_OUT_4 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1632 134 DFF_OUT_1 DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1633 133 DFF_OUT_0 DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1634 VDD 135 132 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1635 VDD 134 131 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1636 VDD 133 130 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1637 126 135 129 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1638 125 134 128 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1639 124 133 127 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=145.799998051317E-15 PD=1.4400000054593E-6 
+PS=539.999973625527E-9 M=1 
M1640 _DFF_OUT_6 _DFF_OUT_5 126 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1641 _DFF_OUT_6 _DFF_OUT_5 125 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1642 _DFF_OUT_6 _DFF_OUT_4 124 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=243.000010304723E-15 AS=145.799998051317E-15 
+PD=1.4400000054593E-6 PS=539.999973625527E-9 M=1 
M1643 127 130 121 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1644 129 132 123 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1645 128 131 122 VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=145.799998051317E-15 PD=539.999973625527E-9 
+PS=539.999973625527E-9 M=1 
M1646 126 DFF_OUT_5 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1647 125 DFF_OUT_5 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1648 124 DFF_OUT_4 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=539.999973625527E-9 AD=145.799998051317E-15 AS=243.000010304723E-15 
+PD=539.999973625527E-9 PS=1.4400000054593E-6 M=1 
M1649 123 126 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1650 122 125 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1651 121 124 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=145.799998051317E-15 AS=243.000010304723E-15 PD=539.999973625527E-9 
+PS=1.4400000054593E-6 M=1 
M1652 120 112 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1653 150 151 H_0 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1654 149 151 H_1 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1655 148 151 H_2 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1656 147 151 H_3 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1657 H_1 142 DFF_OUT_4 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1658 H_1 146 _DFF_OUT_4 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1659 H_2 141 DFF_OUT_5 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1660 H_2 145 _DFF_OUT_5 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1661 H_0 140 DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1662 H_0 144 _DFF_OUT_2 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1663 H_3 139 DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1664 H_3 143 _DFF_OUT_6 VDD  TSMC18DP  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1665 100 111 6 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1666 99 111 90 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1667 98 111 5 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1668 97 111 89 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1669 96 111 4 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1670 95 111 88 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1671 94 111 3 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1672 VDD 109 83 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1673 VDD 109 82 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1674 VDD 109 81 VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1675 13 109 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1676 12 109 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1677 11 109 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1678 10 109 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1679 157 152 153 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1680 160 152 156 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1681 159 152 155 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1682 158 152 154 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1683 117 112 105 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1684 116 112 104 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1685 115 112 103 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1686 114 112 102 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1687 113 112 101 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1688 119 112 107 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1689 118 112 106 VDD  TSMC18DP  L=180.000000682412E-9 W=720.000002729648E-9 
+AD=323.999995669594E-15 AS=323.999995669594E-15 PD=1.62000003456342E-6 
+PS=1.62000003456342E-6 M=1 
M1690 160 164 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1691 159 163 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1692 158 162 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1693 157 161 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1694 119 _DFF_OUT_6 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1695 118 _DFF_OUT_5 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1696 117 _DFF_OUT_4 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1697 116 _DFF_OUT_3 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1698 115 _DFF_OUT_2 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1699 114 _DFF_OUT_1 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1700 113 _DFF_OUT_0 VDD VDD  TSMC18DP  L=360.000001364824E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1701 94 101 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1702 100 107 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1703 99 106 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1704 98 105 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1705 97 104 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1706 96 103 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1707 95 102 VDD VDD  TSMC18DP  L=360.000001364824E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1708 OUT_0 164 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1709 OUT_1 163 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1710 OUT_2 162 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1711 OUT_3 161 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1712 164 160 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1713 163 159 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1714 162 158 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1715 161 157 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1716 156 150 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1717 155 149 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1718 154 148 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1719 153 147 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1720 152 151 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1721 151 120 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1722 90 83 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1723 89 82 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1724 88 81 VDD VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1725 VDD 10 3 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1726 VDD 13 6 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1727 VDD 12 5 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1728 VDD 11 4 VDD  TSMC18DP  L=180.000000682412E-9 W=1.07999994725105E-6 
+AD=486.000020609445E-15 AS=486.000020609445E-15 PD=1.97999997908482E-6 
+PS=1.97999997908482E-6 M=1 
M1729 86 92 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1730 85 91 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1731 65 72 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1732 64 71 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1733 8 15 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1734 7 14 GND GND  TSMC18DN  L=180.000000682412E-9 W=1.62000003456342E-6 
+AD=728.999976704059E-15 AS=728.999976704059E-15 PD=2.51999995271035E-6 
+PS=2.51999995271035E-6 M=1 
M1735 87 86 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1736 66 65 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1737 9 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1738 92 86 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1739 91 85 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1740 72 65 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1741 71 64 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1742 15 8 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1743 14 7 GND GND  TSMC18DN  L=1.4400000054593E-6 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1744 109 108 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1745 108 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1746 91 110 A0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1747 71 110 A1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1748 14 110 A2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1749 112 111 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1750 111 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1751 110 CLK GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1752 92 CLK 85 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1753 72 CLK 64 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1754 15 CLK 7 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1755 _DFF_OUT_6 119 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1756 _DFF_OUT_5 118 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1757 _DFF_OUT_4 117 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1758 _DFF_OUT_3 116 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1759 _DFF_OUT_2 115 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1760 _DFF_OUT_1 114 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1761 _DFF_OUT_0 113 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=1.35000004775065E-6 AD=607.499998656752E-15 AS=607.499998656752E-15 
+PD=2.25000007958442E-6 PS=2.25000007958442E-6 M=1 
M1762 DFF_OUT_3 _DFF_OUT_3 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1763 DFF_OUT_2 _DFF_OUT_2 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1764 DFF_OUT_1 _DFF_OUT_1 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1765 DFF_OUT_0 _DFF_OUT_0 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1766 DFF_OUT_6 _DFF_OUT_6 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1767 DFF_OUT_5 _DFF_OUT_5 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1768 DFF_OUT_4 _DFF_OUT_4 GND GND  TSMC18DN  L=180.000000682412E-9 
+W=810.000017281709E-9 AD=364.499988352029E-15 AS=364.499988352029E-15 
+PD=1.70999999227206E-6 PS=1.70999999227206E-6 M=1 
M1769 107 100 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1770 106 99 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1771 105 98 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1772 104 97 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1773 103 96 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1774 102 95 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1775 101 94 GND GND  TSMC18DN  L=180.000000682412E-9 W=810.000017281709E-9 
+AD=364.499988352029E-15 AS=364.499988352029E-15 PD=1.70999999227206E-6 
+PS=1.70999999227206E-6 M=1 
M1776 142 129 189 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1777 141 129 188 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1778 189 127 187 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1779 188 128 186 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1780 140 128 185 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1781 187 138 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1782 186 137 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1783 185 127 184 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1784 184 136 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1785 139 129 183 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1786 183 128 182 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1787 182 127 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1788 93 87 181 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1789 181 66 180 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1790 180 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1791 84 66 179 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1792 179 86 178 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1793 178 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1794 76 87 177 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1795 177 65 176 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1796 176 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1797 70 86 175 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1798 175 65 174 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1799 174 8 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1800 28 9 173 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1801 173 86 172 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1802 172 65 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1803 16 87 171 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1804 171 9 170 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1805 170 65 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1806 2 66 169 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1807 169 9 168 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1808 168 86 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1809 1 87 167 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=405.000008139519E-15 AS=161.999997834797E-15 PD=1.7999999499807E-6 
+PS=360.000001364824E-9 M=1 
M1810 167 66 166 GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=161.999997834797E-15 PD=360.000001364824E-9 
+PS=360.000001364824E-9 M=1 
M1811 166 9 GND GND  TSMC18DN  L=180.000000682412E-9 W=899.999974990351E-9 
+AD=161.999997834797E-15 AS=405.000008139519E-15 PD=360.000001364824E-9 
+PS=1.7999999499807E-6 M=1 
M1812 150 152 H_0 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1813 149 152 H_1 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1814 148 152 H_2 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1815 147 152 H_3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1816 H_1 146 DFF_OUT_4 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1817 H_1 142 _DFF_OUT_4 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1818 H_2 145 DFF_OUT_5 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1819 H_2 141 _DFF_OUT_5 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1820 H_0 144 DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1821 H_0 140 _DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1822 H_3 143 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1823 H_3 139 _DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1824 146 142 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1825 145 141 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1826 144 140 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1827 143 139 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1828 138 128 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1829 137 127 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1830 136 129 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1831 _DFF_OUT_4 DFF_OUT_3 135 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1832 _DFF_OUT_2 DFF_OUT_1 134 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1833 _DFF_OUT_2 DFF_OUT_0 133 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1834 135 _DFF_OUT_3 DFF_OUT_4 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1835 134 _DFF_OUT_1 DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1836 133 _DFF_OUT_0 DFF_OUT_2 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1837 GND 135 132 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1838 GND 134 131 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1839 GND 133 130 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1840 126 132 129 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1841 125 131 128 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1842 124 130 127 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1843 _DFF_OUT_6 DFF_OUT_5 126 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1844 _DFF_OUT_6 DFF_OUT_5 125 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1845 _DFF_OUT_6 DFF_OUT_4 124 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=89.0999988091383E-15 
+PD=1.35000004775065E-6 PS=629.999988177588E-9 M=1 
M1846 127 133 121 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1847 129 135 123 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1848 128 134 122 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1849 126 _DFF_OUT_5 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1850 125 _DFF_OUT_5 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1851 124 _DFF_OUT_4 DFF_OUT_6 GND  TSMC18DN  L=180.000000682412E-9 
+W=269.999986812763E-9 AD=89.0999988091383E-15 AS=153.900004719321E-15 
+PD=629.999988177588E-9 PS=1.35000004775065E-6 M=1 
M1852 123 126 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1853 122 125 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1854 121 124 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1855 120 112 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1856 100 112 6 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1857 99 112 90 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1858 98 112 5 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1859 97 112 89 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1860 96 112 4 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1861 95 112 88 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1862 94 112 3 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1863 83 1 83 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1864 82 1 82 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1865 81 1 81 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=153.900004719321E-15 PD=629.999988177588E-9 
+PS=1.35000004775065E-6 M=1 
M1866 83 2 80 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1867 82 2 79 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1868 81 2 74 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1869 80 16 78 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1870 79 16 77 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1871 74 16 74 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1872 77 28 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1873 74 28 74 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1874 78 28 75 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1875 75 93 73 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1876 68 93 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1877 74 93 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1878 73 84 73 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1879 68 84 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1880 67 84 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1881 73 76 73 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1882 68 76 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1883 67 76 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1884 73 70 69 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1885 68 70 68 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1886 67 70 67 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1887 69 109 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1888 68 109 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1889 67 109 GND GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1890 GND 109 63 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1891 GND 109 62 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1892 GND 109 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1893 GND 109 60 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1894 63 70 61 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1895 62 70 58 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1896 57 70 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1897 60 70 60 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1898 61 76 59 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1899 58 76 58 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1900 57 76 57 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1901 60 76 26 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1902 57 84 24 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1903 26 84 26 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1904 59 84 25 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1905 58 84 27 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1906 25 93 25 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1907 27 93 19 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1908 24 93 24 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1909 26 93 23 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1910 23 28 21 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1911 25 28 22 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1912 19 28 19 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1913 24 28 18 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1914 22 16 20 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1915 19 16 19 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1916 18 16 18 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1917 21 16 17 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1918 20 2 13 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1919 19 2 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1920 18 2 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1921 17 2 10 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=89.0999988091383E-15 AS=89.0999988091383E-15 PD=629.999988177588E-9 
+PS=629.999988177588E-9 M=1 
M1922 13 1 13 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1923 12 1 12 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1924 11 1 11 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1925 10 1 10 GND  TSMC18DN  L=180.000000682412E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=89.0999988091383E-15 PD=1.35000004775065E-6 
+PS=629.999988177588E-9 M=1 
M1926 160 164 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1927 159 163 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1928 158 162 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1929 157 161 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1930 119 _DFF_OUT_6 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1931 118 _DFF_OUT_5 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1932 117 _DFF_OUT_4 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1933 116 _DFF_OUT_3 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1934 115 _DFF_OUT_2 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1935 114 _DFF_OUT_1 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1936 113 _DFF_OUT_0 GND GND  TSMC18DN  L=720.000002729648E-9 
+W=269.999986812763E-9 AD=153.900004719321E-15 AS=153.900004719321E-15 
+PD=1.35000004775065E-6 PS=1.35000004775065E-6 M=1 
M1937 94 101 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1938 100 107 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1939 99 106 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1940 98 105 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1941 97 104 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1942 96 103 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1943 95 102 GND GND  TSMC18DN  L=720.000002729648E-9 W=269.999986812763E-9 
+AD=153.900004719321E-15 AS=153.900004719321E-15 PD=1.35000004775065E-6 
+PS=1.35000004775065E-6 M=1 
M1944 OUT_0 164 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1945 OUT_1 163 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1946 OUT_2 162 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1947 OUT_3 161 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1948 164 160 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1949 163 159 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1950 162 158 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1951 161 157 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1952 157 151 153 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1953 160 151 156 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1954 159 151 155 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1955 158 151 154 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1956 156 150 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1957 155 149 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1958 154 148 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1959 153 147 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1960 152 151 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1961 151 120 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1962 115 111 103 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1963 114 111 102 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1964 113 111 101 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1965 119 111 107 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1966 118 111 106 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1967 117 111 105 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1968 116 111 104 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1969 90 83 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1970 89 82 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1971 88 81 GND GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1972 GND 13 6 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1973 GND 12 5 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1974 GND 11 4 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
M1975 GND 10 3 GND  TSMC18DN  L=180.000000682412E-9 W=539.999973625527E-9 
+AD=243.000010304723E-15 AS=243.000010304723E-15 PD=1.4400000054593E-6 
+PS=1.4400000054593E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS PART1_G1 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc18dN" NMOS 
   
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TRAN  5.00000E-11 1.70000E-08 START=  0.0000    
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
+        DELMAX = 1.00000E-10
.END
